# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vssio_hvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vssio_hvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.525000 25.850000 0.845000 26.170000 ;
      LAYER met4 ;
        RECT 0.525000 25.850000 0.845000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 26.280000 0.845000 26.600000 ;
      LAYER met4 ;
        RECT 0.525000 26.280000 0.845000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 26.710000 0.845000 27.030000 ;
      LAYER met4 ;
        RECT 0.525000 26.710000 0.845000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 27.140000 0.845000 27.460000 ;
      LAYER met4 ;
        RECT 0.525000 27.140000 0.845000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 27.570000 0.845000 27.890000 ;
      LAYER met4 ;
        RECT 0.525000 27.570000 0.845000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 28.000000 0.845000 28.320000 ;
      LAYER met4 ;
        RECT 0.525000 28.000000 0.845000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 28.430000 0.845000 28.750000 ;
      LAYER met4 ;
        RECT 0.525000 28.430000 0.845000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 28.860000 0.845000 29.180000 ;
      LAYER met4 ;
        RECT 0.525000 28.860000 0.845000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 29.290000 0.845000 29.610000 ;
      LAYER met4 ;
        RECT 0.525000 29.290000 0.845000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 29.720000 0.845000 30.040000 ;
      LAYER met4 ;
        RECT 0.525000 29.720000 0.845000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 30.150000 0.845000 30.470000 ;
      LAYER met4 ;
        RECT 0.525000 30.150000 0.845000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 175.935000 13.345000 195.055000 ;
      LAYER met4 ;
        RECT 0.625000 175.935000 13.345000 195.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 195.140000 0.945000 195.460000 ;
      LAYER met4 ;
        RECT 0.625000 195.140000 0.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 195.545000 0.945000 195.865000 ;
      LAYER met4 ;
        RECT 0.625000 195.545000 0.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 195.950000 0.945000 196.270000 ;
      LAYER met4 ;
        RECT 0.625000 195.950000 0.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 196.355000 0.945000 196.675000 ;
      LAYER met4 ;
        RECT 0.625000 196.355000 0.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 196.760000 0.945000 197.080000 ;
      LAYER met4 ;
        RECT 0.625000 196.760000 0.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 197.165000 0.945000 197.485000 ;
      LAYER met4 ;
        RECT 0.625000 197.165000 0.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 197.570000 0.945000 197.890000 ;
      LAYER met4 ;
        RECT 0.625000 197.570000 0.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 197.975000 0.945000 198.295000 ;
      LAYER met4 ;
        RECT 0.625000 197.975000 0.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 198.380000 0.945000 198.700000 ;
      LAYER met4 ;
        RECT 0.625000 198.380000 0.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 198.785000 0.945000 199.105000 ;
      LAYER met4 ;
        RECT 0.625000 198.785000 0.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 199.190000 0.945000 199.510000 ;
      LAYER met4 ;
        RECT 0.625000 199.190000 0.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625000 199.595000 0.945000 199.915000 ;
      LAYER met4 ;
        RECT 0.625000 199.595000 0.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 175.995000 0.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 176.395000 0.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 176.795000 0.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 177.195000 0.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 177.595000 0.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 177.995000 0.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 178.395000 0.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 178.795000 0.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 179.195000 0.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 179.595000 0.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 179.995000 0.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 180.395000 0.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 180.795000 0.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 181.195000 0.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 181.595000 0.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 181.995000 0.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 182.395000 0.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 182.795000 0.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 183.195000 0.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 183.595000 0.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 183.995000 0.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 184.395000 0.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 184.795000 0.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 185.195000 0.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 185.595000 0.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 185.995000 0.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 186.395000 0.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 186.795000 0.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 187.195000 0.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 187.595000 0.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 187.995000 0.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 188.395000 0.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 188.795000 0.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 189.195000 0.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 189.595000 0.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 189.995000 0.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 190.395000 0.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 190.795000 0.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 191.195000 0.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 191.595000 0.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 191.995000 0.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 192.395000 0.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 192.795000 0.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 193.195000 0.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 193.595000 0.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 193.995000 0.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 194.395000 0.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.685000 194.795000 0.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 25.850000 1.255000 26.170000 ;
      LAYER met4 ;
        RECT 0.935000 25.850000 1.255000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 26.280000 1.255000 26.600000 ;
      LAYER met4 ;
        RECT 0.935000 26.280000 1.255000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 26.710000 1.255000 27.030000 ;
      LAYER met4 ;
        RECT 0.935000 26.710000 1.255000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 27.140000 1.255000 27.460000 ;
      LAYER met4 ;
        RECT 0.935000 27.140000 1.255000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 27.570000 1.255000 27.890000 ;
      LAYER met4 ;
        RECT 0.935000 27.570000 1.255000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 28.000000 1.255000 28.320000 ;
      LAYER met4 ;
        RECT 0.935000 28.000000 1.255000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 28.430000 1.255000 28.750000 ;
      LAYER met4 ;
        RECT 0.935000 28.430000 1.255000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 28.860000 1.255000 29.180000 ;
      LAYER met4 ;
        RECT 0.935000 28.860000 1.255000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 29.290000 1.255000 29.610000 ;
      LAYER met4 ;
        RECT 0.935000 29.290000 1.255000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 29.720000 1.255000 30.040000 ;
      LAYER met4 ;
        RECT 0.935000 29.720000 1.255000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 30.150000 1.255000 30.470000 ;
      LAYER met4 ;
        RECT 0.935000 30.150000 1.255000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 195.140000 1.345000 195.460000 ;
      LAYER met4 ;
        RECT 1.025000 195.140000 1.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 195.545000 1.345000 195.865000 ;
      LAYER met4 ;
        RECT 1.025000 195.545000 1.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 195.950000 1.345000 196.270000 ;
      LAYER met4 ;
        RECT 1.025000 195.950000 1.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 196.355000 1.345000 196.675000 ;
      LAYER met4 ;
        RECT 1.025000 196.355000 1.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 196.760000 1.345000 197.080000 ;
      LAYER met4 ;
        RECT 1.025000 196.760000 1.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 197.165000 1.345000 197.485000 ;
      LAYER met4 ;
        RECT 1.025000 197.165000 1.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 197.570000 1.345000 197.890000 ;
      LAYER met4 ;
        RECT 1.025000 197.570000 1.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 197.975000 1.345000 198.295000 ;
      LAYER met4 ;
        RECT 1.025000 197.975000 1.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 198.380000 1.345000 198.700000 ;
      LAYER met4 ;
        RECT 1.025000 198.380000 1.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 198.785000 1.345000 199.105000 ;
      LAYER met4 ;
        RECT 1.025000 198.785000 1.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 199.190000 1.345000 199.510000 ;
      LAYER met4 ;
        RECT 1.025000 199.190000 1.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025000 199.595000 1.345000 199.915000 ;
      LAYER met4 ;
        RECT 1.025000 199.595000 1.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 175.995000 1.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 176.395000 1.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 176.795000 1.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 177.195000 1.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 177.595000 1.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 177.995000 1.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 178.395000 1.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 178.795000 1.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 179.195000 1.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 179.595000 1.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 179.995000 1.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 180.395000 1.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 180.795000 1.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 181.195000 1.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 181.595000 1.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 181.995000 1.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 182.395000 1.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 182.795000 1.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 183.195000 1.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 183.595000 1.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 183.995000 1.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 184.395000 1.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 184.795000 1.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 185.195000 1.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 185.595000 1.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 185.995000 1.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 186.395000 1.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 186.795000 1.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 187.195000 1.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 187.595000 1.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 187.995000 1.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 188.395000 1.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 188.795000 1.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 189.195000 1.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 189.595000 1.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 189.995000 1.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 190.395000 1.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 190.795000 1.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 191.195000 1.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 191.595000 1.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 191.995000 1.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 192.395000 1.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 192.795000 1.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 193.195000 1.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 193.595000 1.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 193.995000 1.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 194.395000 1.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 194.795000 1.285000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 25.850000 1.665000 26.170000 ;
      LAYER met4 ;
        RECT 1.345000 25.850000 1.665000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 26.280000 1.665000 26.600000 ;
      LAYER met4 ;
        RECT 1.345000 26.280000 1.665000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 26.710000 1.665000 27.030000 ;
      LAYER met4 ;
        RECT 1.345000 26.710000 1.665000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 27.140000 1.665000 27.460000 ;
      LAYER met4 ;
        RECT 1.345000 27.140000 1.665000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 27.570000 1.665000 27.890000 ;
      LAYER met4 ;
        RECT 1.345000 27.570000 1.665000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 28.000000 1.665000 28.320000 ;
      LAYER met4 ;
        RECT 1.345000 28.000000 1.665000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 28.430000 1.665000 28.750000 ;
      LAYER met4 ;
        RECT 1.345000 28.430000 1.665000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 28.860000 1.665000 29.180000 ;
      LAYER met4 ;
        RECT 1.345000 28.860000 1.665000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 29.290000 1.665000 29.610000 ;
      LAYER met4 ;
        RECT 1.345000 29.290000 1.665000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 29.720000 1.665000 30.040000 ;
      LAYER met4 ;
        RECT 1.345000 29.720000 1.665000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 30.150000 1.665000 30.470000 ;
      LAYER met4 ;
        RECT 1.345000 30.150000 1.665000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 195.140000 1.745000 195.460000 ;
      LAYER met4 ;
        RECT 1.425000 195.140000 1.745000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 195.545000 1.745000 195.865000 ;
      LAYER met4 ;
        RECT 1.425000 195.545000 1.745000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 195.950000 1.745000 196.270000 ;
      LAYER met4 ;
        RECT 1.425000 195.950000 1.745000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 196.355000 1.745000 196.675000 ;
      LAYER met4 ;
        RECT 1.425000 196.355000 1.745000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 196.760000 1.745000 197.080000 ;
      LAYER met4 ;
        RECT 1.425000 196.760000 1.745000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 197.165000 1.745000 197.485000 ;
      LAYER met4 ;
        RECT 1.425000 197.165000 1.745000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 197.570000 1.745000 197.890000 ;
      LAYER met4 ;
        RECT 1.425000 197.570000 1.745000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 197.975000 1.745000 198.295000 ;
      LAYER met4 ;
        RECT 1.425000 197.975000 1.745000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 198.380000 1.745000 198.700000 ;
      LAYER met4 ;
        RECT 1.425000 198.380000 1.745000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 198.785000 1.745000 199.105000 ;
      LAYER met4 ;
        RECT 1.425000 198.785000 1.745000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 199.190000 1.745000 199.510000 ;
      LAYER met4 ;
        RECT 1.425000 199.190000 1.745000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425000 199.595000 1.745000 199.915000 ;
      LAYER met4 ;
        RECT 1.425000 199.595000 1.745000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 175.995000 1.685000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 176.395000 1.685000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 176.795000 1.685000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 177.195000 1.685000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 177.595000 1.685000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 177.995000 1.685000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 178.395000 1.685000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 178.795000 1.685000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 179.195000 1.685000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 179.595000 1.685000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 179.995000 1.685000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 180.395000 1.685000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 180.795000 1.685000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 181.195000 1.685000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 181.595000 1.685000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 181.995000 1.685000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 182.395000 1.685000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 182.795000 1.685000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 183.195000 1.685000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 183.595000 1.685000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 183.995000 1.685000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 184.395000 1.685000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 184.795000 1.685000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 185.195000 1.685000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 185.595000 1.685000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 185.995000 1.685000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 186.395000 1.685000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 186.795000 1.685000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 187.195000 1.685000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 187.595000 1.685000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 187.995000 1.685000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 188.395000 1.685000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 188.795000 1.685000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 189.195000 1.685000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 189.595000 1.685000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 189.995000 1.685000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 190.395000 1.685000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 190.795000 1.685000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 191.195000 1.685000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 191.595000 1.685000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 191.995000 1.685000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 192.395000 1.685000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 192.795000 1.685000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 193.195000 1.685000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 193.595000 1.685000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 193.995000 1.685000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 194.395000 1.685000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.485000 194.795000 1.685000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 25.850000 2.075000 26.170000 ;
      LAYER met4 ;
        RECT 1.755000 25.850000 2.075000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 26.280000 2.075000 26.600000 ;
      LAYER met4 ;
        RECT 1.755000 26.280000 2.075000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 26.710000 2.075000 27.030000 ;
      LAYER met4 ;
        RECT 1.755000 26.710000 2.075000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 27.140000 2.075000 27.460000 ;
      LAYER met4 ;
        RECT 1.755000 27.140000 2.075000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 27.570000 2.075000 27.890000 ;
      LAYER met4 ;
        RECT 1.755000 27.570000 2.075000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 28.000000 2.075000 28.320000 ;
      LAYER met4 ;
        RECT 1.755000 28.000000 2.075000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 28.430000 2.075000 28.750000 ;
      LAYER met4 ;
        RECT 1.755000 28.430000 2.075000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 28.860000 2.075000 29.180000 ;
      LAYER met4 ;
        RECT 1.755000 28.860000 2.075000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 29.290000 2.075000 29.610000 ;
      LAYER met4 ;
        RECT 1.755000 29.290000 2.075000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 29.720000 2.075000 30.040000 ;
      LAYER met4 ;
        RECT 1.755000 29.720000 2.075000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 30.150000 2.075000 30.470000 ;
      LAYER met4 ;
        RECT 1.755000 30.150000 2.075000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 195.140000 2.145000 195.460000 ;
      LAYER met4 ;
        RECT 1.825000 195.140000 2.145000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 195.545000 2.145000 195.865000 ;
      LAYER met4 ;
        RECT 1.825000 195.545000 2.145000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 195.950000 2.145000 196.270000 ;
      LAYER met4 ;
        RECT 1.825000 195.950000 2.145000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 196.355000 2.145000 196.675000 ;
      LAYER met4 ;
        RECT 1.825000 196.355000 2.145000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 196.760000 2.145000 197.080000 ;
      LAYER met4 ;
        RECT 1.825000 196.760000 2.145000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 197.165000 2.145000 197.485000 ;
      LAYER met4 ;
        RECT 1.825000 197.165000 2.145000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 197.570000 2.145000 197.890000 ;
      LAYER met4 ;
        RECT 1.825000 197.570000 2.145000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 197.975000 2.145000 198.295000 ;
      LAYER met4 ;
        RECT 1.825000 197.975000 2.145000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 198.380000 2.145000 198.700000 ;
      LAYER met4 ;
        RECT 1.825000 198.380000 2.145000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 198.785000 2.145000 199.105000 ;
      LAYER met4 ;
        RECT 1.825000 198.785000 2.145000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 199.190000 2.145000 199.510000 ;
      LAYER met4 ;
        RECT 1.825000 199.190000 2.145000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825000 199.595000 2.145000 199.915000 ;
      LAYER met4 ;
        RECT 1.825000 199.595000 2.145000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 175.995000 2.085000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 176.395000 2.085000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 176.795000 2.085000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 177.195000 2.085000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 177.595000 2.085000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 177.995000 2.085000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 178.395000 2.085000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 178.795000 2.085000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 179.195000 2.085000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 179.595000 2.085000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 179.995000 2.085000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 180.395000 2.085000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 180.795000 2.085000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 181.195000 2.085000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 181.595000 2.085000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 181.995000 2.085000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 182.395000 2.085000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 182.795000 2.085000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 183.195000 2.085000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 183.595000 2.085000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 183.995000 2.085000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 184.395000 2.085000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 184.795000 2.085000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 185.195000 2.085000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 185.595000 2.085000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 185.995000 2.085000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 186.395000 2.085000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 186.795000 2.085000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 187.195000 2.085000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 187.595000 2.085000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 187.995000 2.085000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 188.395000 2.085000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 188.795000 2.085000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 189.195000 2.085000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 189.595000 2.085000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 189.995000 2.085000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 190.395000 2.085000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 190.795000 2.085000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 191.195000 2.085000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 191.595000 2.085000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 191.995000 2.085000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 192.395000 2.085000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 192.795000 2.085000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 193.195000 2.085000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 193.595000 2.085000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 193.995000 2.085000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 194.395000 2.085000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885000 194.795000 2.085000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 195.140000 10.545000 195.460000 ;
      LAYER met4 ;
        RECT 10.225000 195.140000 10.545000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 195.545000 10.545000 195.865000 ;
      LAYER met4 ;
        RECT 10.225000 195.545000 10.545000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 195.950000 10.545000 196.270000 ;
      LAYER met4 ;
        RECT 10.225000 195.950000 10.545000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 196.355000 10.545000 196.675000 ;
      LAYER met4 ;
        RECT 10.225000 196.355000 10.545000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 196.760000 10.545000 197.080000 ;
      LAYER met4 ;
        RECT 10.225000 196.760000 10.545000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 197.165000 10.545000 197.485000 ;
      LAYER met4 ;
        RECT 10.225000 197.165000 10.545000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 197.570000 10.545000 197.890000 ;
      LAYER met4 ;
        RECT 10.225000 197.570000 10.545000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 197.975000 10.545000 198.295000 ;
      LAYER met4 ;
        RECT 10.225000 197.975000 10.545000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 198.380000 10.545000 198.700000 ;
      LAYER met4 ;
        RECT 10.225000 198.380000 10.545000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 198.785000 10.545000 199.105000 ;
      LAYER met4 ;
        RECT 10.225000 198.785000 10.545000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 199.190000 10.545000 199.510000 ;
      LAYER met4 ;
        RECT 10.225000 199.190000 10.545000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225000 199.595000 10.545000 199.915000 ;
      LAYER met4 ;
        RECT 10.225000 199.595000 10.545000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 25.850000 10.595000 26.170000 ;
      LAYER met4 ;
        RECT 10.275000 25.850000 10.595000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 26.280000 10.595000 26.600000 ;
      LAYER met4 ;
        RECT 10.275000 26.280000 10.595000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 26.710000 10.595000 27.030000 ;
      LAYER met4 ;
        RECT 10.275000 26.710000 10.595000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 27.140000 10.595000 27.460000 ;
      LAYER met4 ;
        RECT 10.275000 27.140000 10.595000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 27.570000 10.595000 27.890000 ;
      LAYER met4 ;
        RECT 10.275000 27.570000 10.595000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 28.000000 10.595000 28.320000 ;
      LAYER met4 ;
        RECT 10.275000 28.000000 10.595000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 28.430000 10.595000 28.750000 ;
      LAYER met4 ;
        RECT 10.275000 28.430000 10.595000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 28.860000 10.595000 29.180000 ;
      LAYER met4 ;
        RECT 10.275000 28.860000 10.595000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 29.290000 10.595000 29.610000 ;
      LAYER met4 ;
        RECT 10.275000 29.290000 10.595000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 29.720000 10.595000 30.040000 ;
      LAYER met4 ;
        RECT 10.275000 29.720000 10.595000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 30.150000 10.595000 30.470000 ;
      LAYER met4 ;
        RECT 10.275000 30.150000 10.595000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 175.995000 10.485000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 176.395000 10.485000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 176.795000 10.485000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 177.195000 10.485000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 177.595000 10.485000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 177.995000 10.485000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 178.395000 10.485000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 178.795000 10.485000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 179.195000 10.485000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 179.595000 10.485000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 179.995000 10.485000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 180.395000 10.485000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 180.795000 10.485000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 181.195000 10.485000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 181.595000 10.485000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 181.995000 10.485000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 182.395000 10.485000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 182.795000 10.485000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 183.195000 10.485000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 183.595000 10.485000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 183.995000 10.485000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 184.395000 10.485000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 184.795000 10.485000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 185.195000 10.485000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 185.595000 10.485000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 185.995000 10.485000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 186.395000 10.485000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 186.795000 10.485000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 187.195000 10.485000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 187.595000 10.485000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 187.995000 10.485000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 188.395000 10.485000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 188.795000 10.485000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 189.195000 10.485000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 189.595000 10.485000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 189.995000 10.485000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 190.395000 10.485000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 190.795000 10.485000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 191.195000 10.485000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 191.595000 10.485000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 191.995000 10.485000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 192.395000 10.485000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 192.795000 10.485000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 193.195000 10.485000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 193.595000 10.485000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 193.995000 10.485000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 194.395000 10.485000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.285000 194.795000 10.485000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 195.140000 10.945000 195.460000 ;
      LAYER met4 ;
        RECT 10.625000 195.140000 10.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 195.545000 10.945000 195.865000 ;
      LAYER met4 ;
        RECT 10.625000 195.545000 10.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 195.950000 10.945000 196.270000 ;
      LAYER met4 ;
        RECT 10.625000 195.950000 10.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 196.355000 10.945000 196.675000 ;
      LAYER met4 ;
        RECT 10.625000 196.355000 10.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 196.760000 10.945000 197.080000 ;
      LAYER met4 ;
        RECT 10.625000 196.760000 10.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 197.165000 10.945000 197.485000 ;
      LAYER met4 ;
        RECT 10.625000 197.165000 10.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 197.570000 10.945000 197.890000 ;
      LAYER met4 ;
        RECT 10.625000 197.570000 10.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 197.975000 10.945000 198.295000 ;
      LAYER met4 ;
        RECT 10.625000 197.975000 10.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 198.380000 10.945000 198.700000 ;
      LAYER met4 ;
        RECT 10.625000 198.380000 10.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 198.785000 10.945000 199.105000 ;
      LAYER met4 ;
        RECT 10.625000 198.785000 10.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 199.190000 10.945000 199.510000 ;
      LAYER met4 ;
        RECT 10.625000 199.190000 10.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625000 199.595000 10.945000 199.915000 ;
      LAYER met4 ;
        RECT 10.625000 199.595000 10.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 25.850000 11.000000 26.170000 ;
      LAYER met4 ;
        RECT 10.680000 25.850000 11.000000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 26.280000 11.000000 26.600000 ;
      LAYER met4 ;
        RECT 10.680000 26.280000 11.000000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 26.710000 11.000000 27.030000 ;
      LAYER met4 ;
        RECT 10.680000 26.710000 11.000000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 27.140000 11.000000 27.460000 ;
      LAYER met4 ;
        RECT 10.680000 27.140000 11.000000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 27.570000 11.000000 27.890000 ;
      LAYER met4 ;
        RECT 10.680000 27.570000 11.000000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 28.000000 11.000000 28.320000 ;
      LAYER met4 ;
        RECT 10.680000 28.000000 11.000000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 28.430000 11.000000 28.750000 ;
      LAYER met4 ;
        RECT 10.680000 28.430000 11.000000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 28.860000 11.000000 29.180000 ;
      LAYER met4 ;
        RECT 10.680000 28.860000 11.000000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 29.290000 11.000000 29.610000 ;
      LAYER met4 ;
        RECT 10.680000 29.290000 11.000000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 29.720000 11.000000 30.040000 ;
      LAYER met4 ;
        RECT 10.680000 29.720000 11.000000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 30.150000 11.000000 30.470000 ;
      LAYER met4 ;
        RECT 10.680000 30.150000 11.000000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 175.995000 10.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 176.395000 10.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 176.795000 10.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 177.195000 10.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 177.595000 10.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 177.995000 10.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 178.395000 10.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 178.795000 10.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 179.195000 10.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 179.595000 10.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 179.995000 10.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 180.395000 10.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 180.795000 10.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 181.195000 10.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 181.595000 10.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 181.995000 10.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 182.395000 10.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 182.795000 10.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 183.195000 10.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 183.595000 10.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 183.995000 10.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 184.395000 10.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 184.795000 10.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 185.195000 10.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 185.595000 10.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 185.995000 10.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 186.395000 10.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 186.795000 10.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 187.195000 10.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 187.595000 10.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 187.995000 10.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 188.395000 10.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 188.795000 10.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 189.195000 10.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 189.595000 10.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 189.995000 10.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 190.395000 10.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 190.795000 10.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 191.195000 10.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 191.595000 10.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 191.995000 10.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 192.395000 10.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 192.795000 10.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 193.195000 10.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 193.595000 10.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 193.995000 10.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 194.395000 10.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 194.795000 10.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 195.140000 11.345000 195.460000 ;
      LAYER met4 ;
        RECT 11.025000 195.140000 11.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 195.545000 11.345000 195.865000 ;
      LAYER met4 ;
        RECT 11.025000 195.545000 11.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 195.950000 11.345000 196.270000 ;
      LAYER met4 ;
        RECT 11.025000 195.950000 11.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 196.355000 11.345000 196.675000 ;
      LAYER met4 ;
        RECT 11.025000 196.355000 11.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 196.760000 11.345000 197.080000 ;
      LAYER met4 ;
        RECT 11.025000 196.760000 11.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 197.165000 11.345000 197.485000 ;
      LAYER met4 ;
        RECT 11.025000 197.165000 11.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 197.570000 11.345000 197.890000 ;
      LAYER met4 ;
        RECT 11.025000 197.570000 11.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 197.975000 11.345000 198.295000 ;
      LAYER met4 ;
        RECT 11.025000 197.975000 11.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 198.380000 11.345000 198.700000 ;
      LAYER met4 ;
        RECT 11.025000 198.380000 11.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 198.785000 11.345000 199.105000 ;
      LAYER met4 ;
        RECT 11.025000 198.785000 11.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 199.190000 11.345000 199.510000 ;
      LAYER met4 ;
        RECT 11.025000 199.190000 11.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025000 199.595000 11.345000 199.915000 ;
      LAYER met4 ;
        RECT 11.025000 199.595000 11.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 175.995000 11.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 176.395000 11.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 176.795000 11.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 177.195000 11.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 177.595000 11.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 177.995000 11.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 178.395000 11.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 178.795000 11.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 179.195000 11.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 179.595000 11.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 179.995000 11.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 180.395000 11.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 180.795000 11.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 181.195000 11.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 181.595000 11.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 181.995000 11.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 182.395000 11.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 182.795000 11.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 183.195000 11.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 183.595000 11.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 183.995000 11.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 184.395000 11.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 184.795000 11.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 185.195000 11.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 185.595000 11.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 185.995000 11.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 186.395000 11.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 186.795000 11.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 187.195000 11.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 187.595000 11.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 187.995000 11.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 188.395000 11.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 188.795000 11.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 189.195000 11.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 189.595000 11.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 189.995000 11.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 190.395000 11.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 190.795000 11.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 191.195000 11.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 191.595000 11.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 191.995000 11.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 192.395000 11.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 192.795000 11.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 193.195000 11.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 193.595000 11.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 193.995000 11.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 194.395000 11.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 194.795000 11.285000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 25.850000 11.405000 26.170000 ;
      LAYER met4 ;
        RECT 11.085000 25.850000 11.405000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 26.280000 11.405000 26.600000 ;
      LAYER met4 ;
        RECT 11.085000 26.280000 11.405000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 26.710000 11.405000 27.030000 ;
      LAYER met4 ;
        RECT 11.085000 26.710000 11.405000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 27.140000 11.405000 27.460000 ;
      LAYER met4 ;
        RECT 11.085000 27.140000 11.405000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 27.570000 11.405000 27.890000 ;
      LAYER met4 ;
        RECT 11.085000 27.570000 11.405000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 28.000000 11.405000 28.320000 ;
      LAYER met4 ;
        RECT 11.085000 28.000000 11.405000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 28.430000 11.405000 28.750000 ;
      LAYER met4 ;
        RECT 11.085000 28.430000 11.405000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 28.860000 11.405000 29.180000 ;
      LAYER met4 ;
        RECT 11.085000 28.860000 11.405000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 29.290000 11.405000 29.610000 ;
      LAYER met4 ;
        RECT 11.085000 29.290000 11.405000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 29.720000 11.405000 30.040000 ;
      LAYER met4 ;
        RECT 11.085000 29.720000 11.405000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 30.150000 11.405000 30.470000 ;
      LAYER met4 ;
        RECT 11.085000 30.150000 11.405000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 195.140000 11.745000 195.460000 ;
      LAYER met4 ;
        RECT 11.425000 195.140000 11.745000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 195.545000 11.745000 195.865000 ;
      LAYER met4 ;
        RECT 11.425000 195.545000 11.745000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 195.950000 11.745000 196.270000 ;
      LAYER met4 ;
        RECT 11.425000 195.950000 11.745000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 196.355000 11.745000 196.675000 ;
      LAYER met4 ;
        RECT 11.425000 196.355000 11.745000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 196.760000 11.745000 197.080000 ;
      LAYER met4 ;
        RECT 11.425000 196.760000 11.745000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 197.165000 11.745000 197.485000 ;
      LAYER met4 ;
        RECT 11.425000 197.165000 11.745000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 197.570000 11.745000 197.890000 ;
      LAYER met4 ;
        RECT 11.425000 197.570000 11.745000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 197.975000 11.745000 198.295000 ;
      LAYER met4 ;
        RECT 11.425000 197.975000 11.745000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 198.380000 11.745000 198.700000 ;
      LAYER met4 ;
        RECT 11.425000 198.380000 11.745000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 198.785000 11.745000 199.105000 ;
      LAYER met4 ;
        RECT 11.425000 198.785000 11.745000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 199.190000 11.745000 199.510000 ;
      LAYER met4 ;
        RECT 11.425000 199.190000 11.745000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425000 199.595000 11.745000 199.915000 ;
      LAYER met4 ;
        RECT 11.425000 199.595000 11.745000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 175.995000 11.685000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 176.395000 11.685000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 176.795000 11.685000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 177.195000 11.685000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 177.595000 11.685000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 177.995000 11.685000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 178.395000 11.685000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 178.795000 11.685000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 179.195000 11.685000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 179.595000 11.685000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 179.995000 11.685000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 180.395000 11.685000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 180.795000 11.685000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 181.195000 11.685000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 181.595000 11.685000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 181.995000 11.685000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 182.395000 11.685000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 182.795000 11.685000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 183.195000 11.685000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 183.595000 11.685000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 183.995000 11.685000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 184.395000 11.685000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 184.795000 11.685000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 185.195000 11.685000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 185.595000 11.685000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 185.995000 11.685000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 186.395000 11.685000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 186.795000 11.685000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 187.195000 11.685000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 187.595000 11.685000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 187.995000 11.685000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 188.395000 11.685000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 188.795000 11.685000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 189.195000 11.685000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 189.595000 11.685000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 189.995000 11.685000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 190.395000 11.685000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 190.795000 11.685000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 191.195000 11.685000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 191.595000 11.685000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 191.995000 11.685000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 192.395000 11.685000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 192.795000 11.685000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 193.195000 11.685000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 193.595000 11.685000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 193.995000 11.685000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 194.395000 11.685000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.485000 194.795000 11.685000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 25.850000 11.810000 26.170000 ;
      LAYER met4 ;
        RECT 11.490000 25.850000 11.810000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 26.280000 11.810000 26.600000 ;
      LAYER met4 ;
        RECT 11.490000 26.280000 11.810000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 26.710000 11.810000 27.030000 ;
      LAYER met4 ;
        RECT 11.490000 26.710000 11.810000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 27.140000 11.810000 27.460000 ;
      LAYER met4 ;
        RECT 11.490000 27.140000 11.810000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 27.570000 11.810000 27.890000 ;
      LAYER met4 ;
        RECT 11.490000 27.570000 11.810000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 28.000000 11.810000 28.320000 ;
      LAYER met4 ;
        RECT 11.490000 28.000000 11.810000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 28.430000 11.810000 28.750000 ;
      LAYER met4 ;
        RECT 11.490000 28.430000 11.810000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 28.860000 11.810000 29.180000 ;
      LAYER met4 ;
        RECT 11.490000 28.860000 11.810000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 29.290000 11.810000 29.610000 ;
      LAYER met4 ;
        RECT 11.490000 29.290000 11.810000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 29.720000 11.810000 30.040000 ;
      LAYER met4 ;
        RECT 11.490000 29.720000 11.810000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 30.150000 11.810000 30.470000 ;
      LAYER met4 ;
        RECT 11.490000 30.150000 11.810000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 195.140000 12.145000 195.460000 ;
      LAYER met4 ;
        RECT 11.825000 195.140000 12.145000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 195.545000 12.145000 195.865000 ;
      LAYER met4 ;
        RECT 11.825000 195.545000 12.145000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 195.950000 12.145000 196.270000 ;
      LAYER met4 ;
        RECT 11.825000 195.950000 12.145000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 196.355000 12.145000 196.675000 ;
      LAYER met4 ;
        RECT 11.825000 196.355000 12.145000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 196.760000 12.145000 197.080000 ;
      LAYER met4 ;
        RECT 11.825000 196.760000 12.145000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 197.165000 12.145000 197.485000 ;
      LAYER met4 ;
        RECT 11.825000 197.165000 12.145000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 197.570000 12.145000 197.890000 ;
      LAYER met4 ;
        RECT 11.825000 197.570000 12.145000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 197.975000 12.145000 198.295000 ;
      LAYER met4 ;
        RECT 11.825000 197.975000 12.145000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 198.380000 12.145000 198.700000 ;
      LAYER met4 ;
        RECT 11.825000 198.380000 12.145000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 198.785000 12.145000 199.105000 ;
      LAYER met4 ;
        RECT 11.825000 198.785000 12.145000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 199.190000 12.145000 199.510000 ;
      LAYER met4 ;
        RECT 11.825000 199.190000 12.145000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825000 199.595000 12.145000 199.915000 ;
      LAYER met4 ;
        RECT 11.825000 199.595000 12.145000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 175.995000 12.085000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 176.395000 12.085000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 176.795000 12.085000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 177.195000 12.085000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 177.595000 12.085000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 177.995000 12.085000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 178.395000 12.085000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 178.795000 12.085000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 179.195000 12.085000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 179.595000 12.085000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 179.995000 12.085000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 180.395000 12.085000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 180.795000 12.085000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 181.195000 12.085000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 181.595000 12.085000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 181.995000 12.085000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 182.395000 12.085000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 182.795000 12.085000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 183.195000 12.085000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 183.595000 12.085000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 183.995000 12.085000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 184.395000 12.085000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 184.795000 12.085000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 185.195000 12.085000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 185.595000 12.085000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 185.995000 12.085000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 186.395000 12.085000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 186.795000 12.085000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 187.195000 12.085000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 187.595000 12.085000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 187.995000 12.085000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 188.395000 12.085000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 188.795000 12.085000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 189.195000 12.085000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 189.595000 12.085000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 189.995000 12.085000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 190.395000 12.085000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 190.795000 12.085000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 191.195000 12.085000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 191.595000 12.085000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 191.995000 12.085000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 192.395000 12.085000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 192.795000 12.085000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 193.195000 12.085000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 193.595000 12.085000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 193.995000 12.085000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 194.395000 12.085000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.885000 194.795000 12.085000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 25.850000 12.215000 26.170000 ;
      LAYER met4 ;
        RECT 11.895000 25.850000 12.215000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 26.280000 12.215000 26.600000 ;
      LAYER met4 ;
        RECT 11.895000 26.280000 12.215000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 26.710000 12.215000 27.030000 ;
      LAYER met4 ;
        RECT 11.895000 26.710000 12.215000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 27.140000 12.215000 27.460000 ;
      LAYER met4 ;
        RECT 11.895000 27.140000 12.215000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 27.570000 12.215000 27.890000 ;
      LAYER met4 ;
        RECT 11.895000 27.570000 12.215000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 28.000000 12.215000 28.320000 ;
      LAYER met4 ;
        RECT 11.895000 28.000000 12.215000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 28.430000 12.215000 28.750000 ;
      LAYER met4 ;
        RECT 11.895000 28.430000 12.215000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 28.860000 12.215000 29.180000 ;
      LAYER met4 ;
        RECT 11.895000 28.860000 12.215000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 29.290000 12.215000 29.610000 ;
      LAYER met4 ;
        RECT 11.895000 29.290000 12.215000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 29.720000 12.215000 30.040000 ;
      LAYER met4 ;
        RECT 11.895000 29.720000 12.215000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 30.150000 12.215000 30.470000 ;
      LAYER met4 ;
        RECT 11.895000 30.150000 12.215000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 195.140000 12.545000 195.460000 ;
      LAYER met4 ;
        RECT 12.225000 195.140000 12.545000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 195.545000 12.545000 195.865000 ;
      LAYER met4 ;
        RECT 12.225000 195.545000 12.545000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 195.950000 12.545000 196.270000 ;
      LAYER met4 ;
        RECT 12.225000 195.950000 12.545000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 196.355000 12.545000 196.675000 ;
      LAYER met4 ;
        RECT 12.225000 196.355000 12.545000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 196.760000 12.545000 197.080000 ;
      LAYER met4 ;
        RECT 12.225000 196.760000 12.545000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 197.165000 12.545000 197.485000 ;
      LAYER met4 ;
        RECT 12.225000 197.165000 12.545000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 197.570000 12.545000 197.890000 ;
      LAYER met4 ;
        RECT 12.225000 197.570000 12.545000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 197.975000 12.545000 198.295000 ;
      LAYER met4 ;
        RECT 12.225000 197.975000 12.545000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 198.380000 12.545000 198.700000 ;
      LAYER met4 ;
        RECT 12.225000 198.380000 12.545000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 198.785000 12.545000 199.105000 ;
      LAYER met4 ;
        RECT 12.225000 198.785000 12.545000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 199.190000 12.545000 199.510000 ;
      LAYER met4 ;
        RECT 12.225000 199.190000 12.545000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225000 199.595000 12.545000 199.915000 ;
      LAYER met4 ;
        RECT 12.225000 199.595000 12.545000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 175.995000 12.485000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 176.395000 12.485000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 176.795000 12.485000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 177.195000 12.485000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 177.595000 12.485000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 177.995000 12.485000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 178.395000 12.485000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 178.795000 12.485000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 179.195000 12.485000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 179.595000 12.485000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 179.995000 12.485000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 180.395000 12.485000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 180.795000 12.485000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 181.195000 12.485000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 181.595000 12.485000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 181.995000 12.485000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 182.395000 12.485000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 182.795000 12.485000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 183.195000 12.485000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 183.595000 12.485000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 183.995000 12.485000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 184.395000 12.485000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 184.795000 12.485000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 185.195000 12.485000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 185.595000 12.485000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 185.995000 12.485000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 186.395000 12.485000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 186.795000 12.485000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 187.195000 12.485000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 187.595000 12.485000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 187.995000 12.485000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 188.395000 12.485000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 188.795000 12.485000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 189.195000 12.485000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 189.595000 12.485000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 189.995000 12.485000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 190.395000 12.485000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 190.795000 12.485000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 191.195000 12.485000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 191.595000 12.485000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 191.995000 12.485000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 192.395000 12.485000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 192.795000 12.485000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 193.195000 12.485000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 193.595000 12.485000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 193.995000 12.485000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 194.395000 12.485000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.285000 194.795000 12.485000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 25.850000 12.620000 26.170000 ;
      LAYER met4 ;
        RECT 12.300000 25.850000 12.620000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 26.280000 12.620000 26.600000 ;
      LAYER met4 ;
        RECT 12.300000 26.280000 12.620000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 26.710000 12.620000 27.030000 ;
      LAYER met4 ;
        RECT 12.300000 26.710000 12.620000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 27.140000 12.620000 27.460000 ;
      LAYER met4 ;
        RECT 12.300000 27.140000 12.620000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 27.570000 12.620000 27.890000 ;
      LAYER met4 ;
        RECT 12.300000 27.570000 12.620000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 28.000000 12.620000 28.320000 ;
      LAYER met4 ;
        RECT 12.300000 28.000000 12.620000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 28.430000 12.620000 28.750000 ;
      LAYER met4 ;
        RECT 12.300000 28.430000 12.620000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 28.860000 12.620000 29.180000 ;
      LAYER met4 ;
        RECT 12.300000 28.860000 12.620000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 29.290000 12.620000 29.610000 ;
      LAYER met4 ;
        RECT 12.300000 29.290000 12.620000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 29.720000 12.620000 30.040000 ;
      LAYER met4 ;
        RECT 12.300000 29.720000 12.620000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 30.150000 12.620000 30.470000 ;
      LAYER met4 ;
        RECT 12.300000 30.150000 12.620000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 195.140000 12.945000 195.460000 ;
      LAYER met4 ;
        RECT 12.625000 195.140000 12.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 195.545000 12.945000 195.865000 ;
      LAYER met4 ;
        RECT 12.625000 195.545000 12.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 195.950000 12.945000 196.270000 ;
      LAYER met4 ;
        RECT 12.625000 195.950000 12.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 196.355000 12.945000 196.675000 ;
      LAYER met4 ;
        RECT 12.625000 196.355000 12.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 196.760000 12.945000 197.080000 ;
      LAYER met4 ;
        RECT 12.625000 196.760000 12.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 197.165000 12.945000 197.485000 ;
      LAYER met4 ;
        RECT 12.625000 197.165000 12.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 197.570000 12.945000 197.890000 ;
      LAYER met4 ;
        RECT 12.625000 197.570000 12.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 197.975000 12.945000 198.295000 ;
      LAYER met4 ;
        RECT 12.625000 197.975000 12.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 198.380000 12.945000 198.700000 ;
      LAYER met4 ;
        RECT 12.625000 198.380000 12.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 198.785000 12.945000 199.105000 ;
      LAYER met4 ;
        RECT 12.625000 198.785000 12.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 199.190000 12.945000 199.510000 ;
      LAYER met4 ;
        RECT 12.625000 199.190000 12.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625000 199.595000 12.945000 199.915000 ;
      LAYER met4 ;
        RECT 12.625000 199.595000 12.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 175.995000 12.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 176.395000 12.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 176.795000 12.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 177.195000 12.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 177.595000 12.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 177.995000 12.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 178.395000 12.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 178.795000 12.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 179.195000 12.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 179.595000 12.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 179.995000 12.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 180.395000 12.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 180.795000 12.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 181.195000 12.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 181.595000 12.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 181.995000 12.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 182.395000 12.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 182.795000 12.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 183.195000 12.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 183.595000 12.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 183.995000 12.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 184.395000 12.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 184.795000 12.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 185.195000 12.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 185.595000 12.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 185.995000 12.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 186.395000 12.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 186.795000 12.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 187.195000 12.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 187.595000 12.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 187.995000 12.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 188.395000 12.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 188.795000 12.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 189.195000 12.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 189.595000 12.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 189.995000 12.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 190.395000 12.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 190.795000 12.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 191.195000 12.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 191.595000 12.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 191.995000 12.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 192.395000 12.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 192.795000 12.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 193.195000 12.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 193.595000 12.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 193.995000 12.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 194.395000 12.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.685000 194.795000 12.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 25.850000 13.025000 26.170000 ;
      LAYER met4 ;
        RECT 12.705000 25.850000 13.025000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 26.280000 13.025000 26.600000 ;
      LAYER met4 ;
        RECT 12.705000 26.280000 13.025000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 26.710000 13.025000 27.030000 ;
      LAYER met4 ;
        RECT 12.705000 26.710000 13.025000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 27.140000 13.025000 27.460000 ;
      LAYER met4 ;
        RECT 12.705000 27.140000 13.025000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 27.570000 13.025000 27.890000 ;
      LAYER met4 ;
        RECT 12.705000 27.570000 13.025000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 28.000000 13.025000 28.320000 ;
      LAYER met4 ;
        RECT 12.705000 28.000000 13.025000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 28.430000 13.025000 28.750000 ;
      LAYER met4 ;
        RECT 12.705000 28.430000 13.025000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 28.860000 13.025000 29.180000 ;
      LAYER met4 ;
        RECT 12.705000 28.860000 13.025000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 29.290000 13.025000 29.610000 ;
      LAYER met4 ;
        RECT 12.705000 29.290000 13.025000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 29.720000 13.025000 30.040000 ;
      LAYER met4 ;
        RECT 12.705000 29.720000 13.025000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 30.150000 13.025000 30.470000 ;
      LAYER met4 ;
        RECT 12.705000 30.150000 13.025000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 195.140000 13.345000 195.460000 ;
      LAYER met4 ;
        RECT 13.025000 195.140000 13.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 195.545000 13.345000 195.865000 ;
      LAYER met4 ;
        RECT 13.025000 195.545000 13.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 195.950000 13.345000 196.270000 ;
      LAYER met4 ;
        RECT 13.025000 195.950000 13.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 196.355000 13.345000 196.675000 ;
      LAYER met4 ;
        RECT 13.025000 196.355000 13.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 196.760000 13.345000 197.080000 ;
      LAYER met4 ;
        RECT 13.025000 196.760000 13.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 197.165000 13.345000 197.485000 ;
      LAYER met4 ;
        RECT 13.025000 197.165000 13.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 197.570000 13.345000 197.890000 ;
      LAYER met4 ;
        RECT 13.025000 197.570000 13.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 197.975000 13.345000 198.295000 ;
      LAYER met4 ;
        RECT 13.025000 197.975000 13.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 198.380000 13.345000 198.700000 ;
      LAYER met4 ;
        RECT 13.025000 198.380000 13.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 198.785000 13.345000 199.105000 ;
      LAYER met4 ;
        RECT 13.025000 198.785000 13.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 199.190000 13.345000 199.510000 ;
      LAYER met4 ;
        RECT 13.025000 199.190000 13.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025000 199.595000 13.345000 199.915000 ;
      LAYER met4 ;
        RECT 13.025000 199.595000 13.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 175.995000 13.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 176.395000 13.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 176.795000 13.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 177.195000 13.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 177.595000 13.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 177.995000 13.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 178.395000 13.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 178.795000 13.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 179.195000 13.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 179.595000 13.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 179.995000 13.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 180.395000 13.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 180.795000 13.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 181.195000 13.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 181.595000 13.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 181.995000 13.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 182.395000 13.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 182.795000 13.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 183.195000 13.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 183.595000 13.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 183.995000 13.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 184.395000 13.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 184.795000 13.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 185.195000 13.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 185.595000 13.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 185.995000 13.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 186.395000 13.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 186.795000 13.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 187.195000 13.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 187.595000 13.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 187.995000 13.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 188.395000 13.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 188.795000 13.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 189.195000 13.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 189.595000 13.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 189.995000 13.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 190.395000 13.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 190.795000 13.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 191.195000 13.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 191.595000 13.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 191.995000 13.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 192.395000 13.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 192.795000 13.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 193.195000 13.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 193.595000 13.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 193.995000 13.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.085000 194.395000 13.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 25.850000 13.430000 26.170000 ;
      LAYER met4 ;
        RECT 13.110000 25.850000 13.430000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 26.280000 13.430000 26.600000 ;
      LAYER met4 ;
        RECT 13.110000 26.280000 13.430000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 26.710000 13.430000 27.030000 ;
      LAYER met4 ;
        RECT 13.110000 26.710000 13.430000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 27.140000 13.430000 27.460000 ;
      LAYER met4 ;
        RECT 13.110000 27.140000 13.430000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 27.570000 13.430000 27.890000 ;
      LAYER met4 ;
        RECT 13.110000 27.570000 13.430000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 28.000000 13.430000 28.320000 ;
      LAYER met4 ;
        RECT 13.110000 28.000000 13.430000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 28.430000 13.430000 28.750000 ;
      LAYER met4 ;
        RECT 13.110000 28.430000 13.430000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 28.860000 13.430000 29.180000 ;
      LAYER met4 ;
        RECT 13.110000 28.860000 13.430000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 29.290000 13.430000 29.610000 ;
      LAYER met4 ;
        RECT 13.110000 29.290000 13.430000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 29.720000 13.430000 30.040000 ;
      LAYER met4 ;
        RECT 13.110000 29.720000 13.430000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 30.150000 13.430000 30.470000 ;
      LAYER met4 ;
        RECT 13.110000 30.150000 13.430000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 25.850000 13.835000 26.170000 ;
      LAYER met4 ;
        RECT 13.515000 25.850000 13.835000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 26.280000 13.835000 26.600000 ;
      LAYER met4 ;
        RECT 13.515000 26.280000 13.835000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 26.710000 13.835000 27.030000 ;
      LAYER met4 ;
        RECT 13.515000 26.710000 13.835000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 27.140000 13.835000 27.460000 ;
      LAYER met4 ;
        RECT 13.515000 27.140000 13.835000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 27.570000 13.835000 27.890000 ;
      LAYER met4 ;
        RECT 13.515000 27.570000 13.835000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 28.000000 13.835000 28.320000 ;
      LAYER met4 ;
        RECT 13.515000 28.000000 13.835000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 28.430000 13.835000 28.750000 ;
      LAYER met4 ;
        RECT 13.515000 28.430000 13.835000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 28.860000 13.835000 29.180000 ;
      LAYER met4 ;
        RECT 13.515000 28.860000 13.835000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 29.290000 13.835000 29.610000 ;
      LAYER met4 ;
        RECT 13.515000 29.290000 13.835000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 29.720000 13.835000 30.040000 ;
      LAYER met4 ;
        RECT 13.515000 29.720000 13.835000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 30.150000 13.835000 30.470000 ;
      LAYER met4 ;
        RECT 13.515000 30.150000 13.835000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 197.190000 13.955000 197.510000 ;
      LAYER met4 ;
        RECT 13.635000 197.190000 13.955000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 197.590000 13.955000 197.910000 ;
      LAYER met4 ;
        RECT 13.635000 197.590000 13.955000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 197.990000 13.955000 198.310000 ;
      LAYER met4 ;
        RECT 13.635000 197.990000 13.955000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 198.390000 13.955000 198.710000 ;
      LAYER met4 ;
        RECT 13.635000 198.390000 13.955000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 198.790000 13.955000 199.110000 ;
      LAYER met4 ;
        RECT 13.635000 198.790000 13.955000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 199.190000 13.955000 199.510000 ;
      LAYER met4 ;
        RECT 13.635000 199.190000 13.955000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635000 199.590000 13.955000 199.910000 ;
      LAYER met4 ;
        RECT 13.635000 199.590000 13.955000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.765000 196.235000 14.085000 196.555000 ;
      LAYER met4 ;
        RECT 13.765000 196.235000 14.085000 196.555000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.765000 196.645000 14.085000 196.965000 ;
      LAYER met4 ;
        RECT 13.765000 196.645000 14.085000 196.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 25.850000 14.240000 26.170000 ;
      LAYER met4 ;
        RECT 13.920000 25.850000 14.240000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 26.280000 14.240000 26.600000 ;
      LAYER met4 ;
        RECT 13.920000 26.280000 14.240000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 26.710000 14.240000 27.030000 ;
      LAYER met4 ;
        RECT 13.920000 26.710000 14.240000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 27.140000 14.240000 27.460000 ;
      LAYER met4 ;
        RECT 13.920000 27.140000 14.240000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 27.570000 14.240000 27.890000 ;
      LAYER met4 ;
        RECT 13.920000 27.570000 14.240000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 28.000000 14.240000 28.320000 ;
      LAYER met4 ;
        RECT 13.920000 28.000000 14.240000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 28.430000 14.240000 28.750000 ;
      LAYER met4 ;
        RECT 13.920000 28.430000 14.240000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 28.860000 14.240000 29.180000 ;
      LAYER met4 ;
        RECT 13.920000 28.860000 14.240000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 29.290000 14.240000 29.610000 ;
      LAYER met4 ;
        RECT 13.920000 29.290000 14.240000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 29.720000 14.240000 30.040000 ;
      LAYER met4 ;
        RECT 13.920000 29.720000 14.240000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 30.150000 14.240000 30.470000 ;
      LAYER met4 ;
        RECT 13.920000 30.150000 14.240000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 197.190000 14.360000 197.510000 ;
      LAYER met4 ;
        RECT 14.040000 197.190000 14.360000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 197.590000 14.360000 197.910000 ;
      LAYER met4 ;
        RECT 14.040000 197.590000 14.360000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 197.990000 14.360000 198.310000 ;
      LAYER met4 ;
        RECT 14.040000 197.990000 14.360000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 198.390000 14.360000 198.710000 ;
      LAYER met4 ;
        RECT 14.040000 198.390000 14.360000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 198.790000 14.360000 199.110000 ;
      LAYER met4 ;
        RECT 14.040000 198.790000 14.360000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 199.190000 14.360000 199.510000 ;
      LAYER met4 ;
        RECT 14.040000 199.190000 14.360000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040000 199.590000 14.360000 199.910000 ;
      LAYER met4 ;
        RECT 14.040000 199.590000 14.360000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 25.850000 14.645000 26.170000 ;
      LAYER met4 ;
        RECT 14.325000 25.850000 14.645000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 26.280000 14.645000 26.600000 ;
      LAYER met4 ;
        RECT 14.325000 26.280000 14.645000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 26.710000 14.645000 27.030000 ;
      LAYER met4 ;
        RECT 14.325000 26.710000 14.645000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 27.140000 14.645000 27.460000 ;
      LAYER met4 ;
        RECT 14.325000 27.140000 14.645000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 27.570000 14.645000 27.890000 ;
      LAYER met4 ;
        RECT 14.325000 27.570000 14.645000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 28.000000 14.645000 28.320000 ;
      LAYER met4 ;
        RECT 14.325000 28.000000 14.645000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 28.430000 14.645000 28.750000 ;
      LAYER met4 ;
        RECT 14.325000 28.430000 14.645000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 28.860000 14.645000 29.180000 ;
      LAYER met4 ;
        RECT 14.325000 28.860000 14.645000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 29.290000 14.645000 29.610000 ;
      LAYER met4 ;
        RECT 14.325000 29.290000 14.645000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 29.720000 14.645000 30.040000 ;
      LAYER met4 ;
        RECT 14.325000 29.720000 14.645000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 30.150000 14.645000 30.470000 ;
      LAYER met4 ;
        RECT 14.325000 30.150000 14.645000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 197.190000 14.765000 197.510000 ;
      LAYER met4 ;
        RECT 14.445000 197.190000 14.765000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 197.590000 14.765000 197.910000 ;
      LAYER met4 ;
        RECT 14.445000 197.590000 14.765000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 197.990000 14.765000 198.310000 ;
      LAYER met4 ;
        RECT 14.445000 197.990000 14.765000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 198.390000 14.765000 198.710000 ;
      LAYER met4 ;
        RECT 14.445000 198.390000 14.765000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 198.790000 14.765000 199.110000 ;
      LAYER met4 ;
        RECT 14.445000 198.790000 14.765000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 199.190000 14.765000 199.510000 ;
      LAYER met4 ;
        RECT 14.445000 199.190000 14.765000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445000 199.590000 14.765000 199.910000 ;
      LAYER met4 ;
        RECT 14.445000 199.590000 14.765000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 25.850000 15.050000 26.170000 ;
      LAYER met4 ;
        RECT 14.730000 25.850000 15.050000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 26.280000 15.050000 26.600000 ;
      LAYER met4 ;
        RECT 14.730000 26.280000 15.050000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 26.710000 15.050000 27.030000 ;
      LAYER met4 ;
        RECT 14.730000 26.710000 15.050000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 27.140000 15.050000 27.460000 ;
      LAYER met4 ;
        RECT 14.730000 27.140000 15.050000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 27.570000 15.050000 27.890000 ;
      LAYER met4 ;
        RECT 14.730000 27.570000 15.050000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 28.000000 15.050000 28.320000 ;
      LAYER met4 ;
        RECT 14.730000 28.000000 15.050000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 28.430000 15.050000 28.750000 ;
      LAYER met4 ;
        RECT 14.730000 28.430000 15.050000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 28.860000 15.050000 29.180000 ;
      LAYER met4 ;
        RECT 14.730000 28.860000 15.050000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 29.290000 15.050000 29.610000 ;
      LAYER met4 ;
        RECT 14.730000 29.290000 15.050000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 29.720000 15.050000 30.040000 ;
      LAYER met4 ;
        RECT 14.730000 29.720000 15.050000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 30.150000 15.050000 30.470000 ;
      LAYER met4 ;
        RECT 14.730000 30.150000 15.050000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 197.190000 15.170000 197.510000 ;
      LAYER met4 ;
        RECT 14.850000 197.190000 15.170000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 197.590000 15.170000 197.910000 ;
      LAYER met4 ;
        RECT 14.850000 197.590000 15.170000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 197.990000 15.170000 198.310000 ;
      LAYER met4 ;
        RECT 14.850000 197.990000 15.170000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 198.390000 15.170000 198.710000 ;
      LAYER met4 ;
        RECT 14.850000 198.390000 15.170000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 198.790000 15.170000 199.110000 ;
      LAYER met4 ;
        RECT 14.850000 198.790000 15.170000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 199.190000 15.170000 199.510000 ;
      LAYER met4 ;
        RECT 14.850000 199.190000 15.170000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850000 199.590000 15.170000 199.910000 ;
      LAYER met4 ;
        RECT 14.850000 199.590000 15.170000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 25.850000 15.455000 26.170000 ;
      LAYER met4 ;
        RECT 15.135000 25.850000 15.455000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 26.280000 15.455000 26.600000 ;
      LAYER met4 ;
        RECT 15.135000 26.280000 15.455000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 26.710000 15.455000 27.030000 ;
      LAYER met4 ;
        RECT 15.135000 26.710000 15.455000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 27.140000 15.455000 27.460000 ;
      LAYER met4 ;
        RECT 15.135000 27.140000 15.455000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 27.570000 15.455000 27.890000 ;
      LAYER met4 ;
        RECT 15.135000 27.570000 15.455000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 28.000000 15.455000 28.320000 ;
      LAYER met4 ;
        RECT 15.135000 28.000000 15.455000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 28.430000 15.455000 28.750000 ;
      LAYER met4 ;
        RECT 15.135000 28.430000 15.455000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 28.860000 15.455000 29.180000 ;
      LAYER met4 ;
        RECT 15.135000 28.860000 15.455000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 29.290000 15.455000 29.610000 ;
      LAYER met4 ;
        RECT 15.135000 29.290000 15.455000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 29.720000 15.455000 30.040000 ;
      LAYER met4 ;
        RECT 15.135000 29.720000 15.455000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 30.150000 15.455000 30.470000 ;
      LAYER met4 ;
        RECT 15.135000 30.150000 15.455000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 197.190000 15.575000 197.510000 ;
      LAYER met4 ;
        RECT 15.255000 197.190000 15.575000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 197.590000 15.575000 197.910000 ;
      LAYER met4 ;
        RECT 15.255000 197.590000 15.575000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 197.990000 15.575000 198.310000 ;
      LAYER met4 ;
        RECT 15.255000 197.990000 15.575000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 198.390000 15.575000 198.710000 ;
      LAYER met4 ;
        RECT 15.255000 198.390000 15.575000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 198.790000 15.575000 199.110000 ;
      LAYER met4 ;
        RECT 15.255000 198.790000 15.575000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 199.190000 15.575000 199.510000 ;
      LAYER met4 ;
        RECT 15.255000 199.190000 15.575000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255000 199.590000 15.575000 199.910000 ;
      LAYER met4 ;
        RECT 15.255000 199.590000 15.575000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 25.850000 15.860000 26.170000 ;
      LAYER met4 ;
        RECT 15.540000 25.850000 15.860000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 26.280000 15.860000 26.600000 ;
      LAYER met4 ;
        RECT 15.540000 26.280000 15.860000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 26.710000 15.860000 27.030000 ;
      LAYER met4 ;
        RECT 15.540000 26.710000 15.860000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 27.140000 15.860000 27.460000 ;
      LAYER met4 ;
        RECT 15.540000 27.140000 15.860000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 27.570000 15.860000 27.890000 ;
      LAYER met4 ;
        RECT 15.540000 27.570000 15.860000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 28.000000 15.860000 28.320000 ;
      LAYER met4 ;
        RECT 15.540000 28.000000 15.860000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 28.430000 15.860000 28.750000 ;
      LAYER met4 ;
        RECT 15.540000 28.430000 15.860000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 28.860000 15.860000 29.180000 ;
      LAYER met4 ;
        RECT 15.540000 28.860000 15.860000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 29.290000 15.860000 29.610000 ;
      LAYER met4 ;
        RECT 15.540000 29.290000 15.860000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 29.720000 15.860000 30.040000 ;
      LAYER met4 ;
        RECT 15.540000 29.720000 15.860000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 30.150000 15.860000 30.470000 ;
      LAYER met4 ;
        RECT 15.540000 30.150000 15.860000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 197.190000 15.980000 197.510000 ;
      LAYER met4 ;
        RECT 15.660000 197.190000 15.980000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 197.590000 15.980000 197.910000 ;
      LAYER met4 ;
        RECT 15.660000 197.590000 15.980000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 197.990000 15.980000 198.310000 ;
      LAYER met4 ;
        RECT 15.660000 197.990000 15.980000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 198.390000 15.980000 198.710000 ;
      LAYER met4 ;
        RECT 15.660000 198.390000 15.980000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 198.790000 15.980000 199.110000 ;
      LAYER met4 ;
        RECT 15.660000 198.790000 15.980000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 199.190000 15.980000 199.510000 ;
      LAYER met4 ;
        RECT 15.660000 199.190000 15.980000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660000 199.590000 15.980000 199.910000 ;
      LAYER met4 ;
        RECT 15.660000 199.590000 15.980000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 25.850000 16.265000 26.170000 ;
      LAYER met4 ;
        RECT 15.945000 25.850000 16.265000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 26.280000 16.265000 26.600000 ;
      LAYER met4 ;
        RECT 15.945000 26.280000 16.265000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 26.710000 16.265000 27.030000 ;
      LAYER met4 ;
        RECT 15.945000 26.710000 16.265000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 27.140000 16.265000 27.460000 ;
      LAYER met4 ;
        RECT 15.945000 27.140000 16.265000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 27.570000 16.265000 27.890000 ;
      LAYER met4 ;
        RECT 15.945000 27.570000 16.265000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 28.000000 16.265000 28.320000 ;
      LAYER met4 ;
        RECT 15.945000 28.000000 16.265000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 28.430000 16.265000 28.750000 ;
      LAYER met4 ;
        RECT 15.945000 28.430000 16.265000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 28.860000 16.265000 29.180000 ;
      LAYER met4 ;
        RECT 15.945000 28.860000 16.265000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 29.290000 16.265000 29.610000 ;
      LAYER met4 ;
        RECT 15.945000 29.290000 16.265000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 29.720000 16.265000 30.040000 ;
      LAYER met4 ;
        RECT 15.945000 29.720000 16.265000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 30.150000 16.265000 30.470000 ;
      LAYER met4 ;
        RECT 15.945000 30.150000 16.265000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 197.190000 16.385000 197.510000 ;
      LAYER met4 ;
        RECT 16.065000 197.190000 16.385000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 197.590000 16.385000 197.910000 ;
      LAYER met4 ;
        RECT 16.065000 197.590000 16.385000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 197.990000 16.385000 198.310000 ;
      LAYER met4 ;
        RECT 16.065000 197.990000 16.385000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 198.390000 16.385000 198.710000 ;
      LAYER met4 ;
        RECT 16.065000 198.390000 16.385000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 198.790000 16.385000 199.110000 ;
      LAYER met4 ;
        RECT 16.065000 198.790000 16.385000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 199.190000 16.385000 199.510000 ;
      LAYER met4 ;
        RECT 16.065000 199.190000 16.385000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065000 199.590000 16.385000 199.910000 ;
      LAYER met4 ;
        RECT 16.065000 199.590000 16.385000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 25.850000 16.670000 26.170000 ;
      LAYER met4 ;
        RECT 16.350000 25.850000 16.670000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 26.280000 16.670000 26.600000 ;
      LAYER met4 ;
        RECT 16.350000 26.280000 16.670000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 26.710000 16.670000 27.030000 ;
      LAYER met4 ;
        RECT 16.350000 26.710000 16.670000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 27.140000 16.670000 27.460000 ;
      LAYER met4 ;
        RECT 16.350000 27.140000 16.670000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 27.570000 16.670000 27.890000 ;
      LAYER met4 ;
        RECT 16.350000 27.570000 16.670000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 28.000000 16.670000 28.320000 ;
      LAYER met4 ;
        RECT 16.350000 28.000000 16.670000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 28.430000 16.670000 28.750000 ;
      LAYER met4 ;
        RECT 16.350000 28.430000 16.670000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 28.860000 16.670000 29.180000 ;
      LAYER met4 ;
        RECT 16.350000 28.860000 16.670000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 29.290000 16.670000 29.610000 ;
      LAYER met4 ;
        RECT 16.350000 29.290000 16.670000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 29.720000 16.670000 30.040000 ;
      LAYER met4 ;
        RECT 16.350000 29.720000 16.670000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 30.150000 16.670000 30.470000 ;
      LAYER met4 ;
        RECT 16.350000 30.150000 16.670000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 197.190000 16.790000 197.510000 ;
      LAYER met4 ;
        RECT 16.470000 197.190000 16.790000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 197.590000 16.790000 197.910000 ;
      LAYER met4 ;
        RECT 16.470000 197.590000 16.790000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 197.990000 16.790000 198.310000 ;
      LAYER met4 ;
        RECT 16.470000 197.990000 16.790000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 198.390000 16.790000 198.710000 ;
      LAYER met4 ;
        RECT 16.470000 198.390000 16.790000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 198.790000 16.790000 199.110000 ;
      LAYER met4 ;
        RECT 16.470000 198.790000 16.790000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 199.190000 16.790000 199.510000 ;
      LAYER met4 ;
        RECT 16.470000 199.190000 16.790000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470000 199.590000 16.790000 199.910000 ;
      LAYER met4 ;
        RECT 16.470000 199.590000 16.790000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 25.850000 17.075000 26.170000 ;
      LAYER met4 ;
        RECT 16.755000 25.850000 17.075000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 26.280000 17.075000 26.600000 ;
      LAYER met4 ;
        RECT 16.755000 26.280000 17.075000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 26.710000 17.075000 27.030000 ;
      LAYER met4 ;
        RECT 16.755000 26.710000 17.075000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 27.140000 17.075000 27.460000 ;
      LAYER met4 ;
        RECT 16.755000 27.140000 17.075000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 27.570000 17.075000 27.890000 ;
      LAYER met4 ;
        RECT 16.755000 27.570000 17.075000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 28.000000 17.075000 28.320000 ;
      LAYER met4 ;
        RECT 16.755000 28.000000 17.075000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 28.430000 17.075000 28.750000 ;
      LAYER met4 ;
        RECT 16.755000 28.430000 17.075000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 28.860000 17.075000 29.180000 ;
      LAYER met4 ;
        RECT 16.755000 28.860000 17.075000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 29.290000 17.075000 29.610000 ;
      LAYER met4 ;
        RECT 16.755000 29.290000 17.075000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 29.720000 17.075000 30.040000 ;
      LAYER met4 ;
        RECT 16.755000 29.720000 17.075000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 30.150000 17.075000 30.470000 ;
      LAYER met4 ;
        RECT 16.755000 30.150000 17.075000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 197.190000 17.195000 197.510000 ;
      LAYER met4 ;
        RECT 16.875000 197.190000 17.195000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 197.590000 17.195000 197.910000 ;
      LAYER met4 ;
        RECT 16.875000 197.590000 17.195000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 197.990000 17.195000 198.310000 ;
      LAYER met4 ;
        RECT 16.875000 197.990000 17.195000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 198.390000 17.195000 198.710000 ;
      LAYER met4 ;
        RECT 16.875000 198.390000 17.195000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 198.790000 17.195000 199.110000 ;
      LAYER met4 ;
        RECT 16.875000 198.790000 17.195000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 199.190000 17.195000 199.510000 ;
      LAYER met4 ;
        RECT 16.875000 199.190000 17.195000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875000 199.590000 17.195000 199.910000 ;
      LAYER met4 ;
        RECT 16.875000 199.590000 17.195000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 25.850000 17.480000 26.170000 ;
      LAYER met4 ;
        RECT 17.160000 25.850000 17.480000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 26.280000 17.480000 26.600000 ;
      LAYER met4 ;
        RECT 17.160000 26.280000 17.480000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 26.710000 17.480000 27.030000 ;
      LAYER met4 ;
        RECT 17.160000 26.710000 17.480000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 27.140000 17.480000 27.460000 ;
      LAYER met4 ;
        RECT 17.160000 27.140000 17.480000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 27.570000 17.480000 27.890000 ;
      LAYER met4 ;
        RECT 17.160000 27.570000 17.480000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 28.000000 17.480000 28.320000 ;
      LAYER met4 ;
        RECT 17.160000 28.000000 17.480000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 28.430000 17.480000 28.750000 ;
      LAYER met4 ;
        RECT 17.160000 28.430000 17.480000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 28.860000 17.480000 29.180000 ;
      LAYER met4 ;
        RECT 17.160000 28.860000 17.480000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 29.290000 17.480000 29.610000 ;
      LAYER met4 ;
        RECT 17.160000 29.290000 17.480000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 29.720000 17.480000 30.040000 ;
      LAYER met4 ;
        RECT 17.160000 29.720000 17.480000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 30.150000 17.480000 30.470000 ;
      LAYER met4 ;
        RECT 17.160000 30.150000 17.480000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 197.190000 17.600000 197.510000 ;
      LAYER met4 ;
        RECT 17.280000 197.190000 17.600000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 197.590000 17.600000 197.910000 ;
      LAYER met4 ;
        RECT 17.280000 197.590000 17.600000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 197.990000 17.600000 198.310000 ;
      LAYER met4 ;
        RECT 17.280000 197.990000 17.600000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 198.390000 17.600000 198.710000 ;
      LAYER met4 ;
        RECT 17.280000 198.390000 17.600000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 198.790000 17.600000 199.110000 ;
      LAYER met4 ;
        RECT 17.280000 198.790000 17.600000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 199.190000 17.600000 199.510000 ;
      LAYER met4 ;
        RECT 17.280000 199.190000 17.600000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280000 199.590000 17.600000 199.910000 ;
      LAYER met4 ;
        RECT 17.280000 199.590000 17.600000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 25.850000 17.885000 26.170000 ;
      LAYER met4 ;
        RECT 17.565000 25.850000 17.885000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 26.280000 17.885000 26.600000 ;
      LAYER met4 ;
        RECT 17.565000 26.280000 17.885000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 26.710000 17.885000 27.030000 ;
      LAYER met4 ;
        RECT 17.565000 26.710000 17.885000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 27.140000 17.885000 27.460000 ;
      LAYER met4 ;
        RECT 17.565000 27.140000 17.885000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 27.570000 17.885000 27.890000 ;
      LAYER met4 ;
        RECT 17.565000 27.570000 17.885000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 28.000000 17.885000 28.320000 ;
      LAYER met4 ;
        RECT 17.565000 28.000000 17.885000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 28.430000 17.885000 28.750000 ;
      LAYER met4 ;
        RECT 17.565000 28.430000 17.885000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 28.860000 17.885000 29.180000 ;
      LAYER met4 ;
        RECT 17.565000 28.860000 17.885000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 29.290000 17.885000 29.610000 ;
      LAYER met4 ;
        RECT 17.565000 29.290000 17.885000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 29.720000 17.885000 30.040000 ;
      LAYER met4 ;
        RECT 17.565000 29.720000 17.885000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 30.150000 17.885000 30.470000 ;
      LAYER met4 ;
        RECT 17.565000 30.150000 17.885000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 197.190000 18.005000 197.510000 ;
      LAYER met4 ;
        RECT 17.685000 197.190000 18.005000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 197.590000 18.005000 197.910000 ;
      LAYER met4 ;
        RECT 17.685000 197.590000 18.005000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 197.990000 18.005000 198.310000 ;
      LAYER met4 ;
        RECT 17.685000 197.990000 18.005000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 198.390000 18.005000 198.710000 ;
      LAYER met4 ;
        RECT 17.685000 198.390000 18.005000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 198.790000 18.005000 199.110000 ;
      LAYER met4 ;
        RECT 17.685000 198.790000 18.005000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 199.190000 18.005000 199.510000 ;
      LAYER met4 ;
        RECT 17.685000 199.190000 18.005000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 199.590000 18.005000 199.910000 ;
      LAYER met4 ;
        RECT 17.685000 199.590000 18.005000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 25.850000 18.290000 26.170000 ;
      LAYER met4 ;
        RECT 17.970000 25.850000 18.290000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 26.280000 18.290000 26.600000 ;
      LAYER met4 ;
        RECT 17.970000 26.280000 18.290000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 26.710000 18.290000 27.030000 ;
      LAYER met4 ;
        RECT 17.970000 26.710000 18.290000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 27.140000 18.290000 27.460000 ;
      LAYER met4 ;
        RECT 17.970000 27.140000 18.290000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 27.570000 18.290000 27.890000 ;
      LAYER met4 ;
        RECT 17.970000 27.570000 18.290000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 28.000000 18.290000 28.320000 ;
      LAYER met4 ;
        RECT 17.970000 28.000000 18.290000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 28.430000 18.290000 28.750000 ;
      LAYER met4 ;
        RECT 17.970000 28.430000 18.290000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 28.860000 18.290000 29.180000 ;
      LAYER met4 ;
        RECT 17.970000 28.860000 18.290000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 29.290000 18.290000 29.610000 ;
      LAYER met4 ;
        RECT 17.970000 29.290000 18.290000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 29.720000 18.290000 30.040000 ;
      LAYER met4 ;
        RECT 17.970000 29.720000 18.290000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 30.150000 18.290000 30.470000 ;
      LAYER met4 ;
        RECT 17.970000 30.150000 18.290000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 197.190000 18.410000 197.510000 ;
      LAYER met4 ;
        RECT 18.090000 197.190000 18.410000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 197.590000 18.410000 197.910000 ;
      LAYER met4 ;
        RECT 18.090000 197.590000 18.410000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 197.990000 18.410000 198.310000 ;
      LAYER met4 ;
        RECT 18.090000 197.990000 18.410000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 198.390000 18.410000 198.710000 ;
      LAYER met4 ;
        RECT 18.090000 198.390000 18.410000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 198.790000 18.410000 199.110000 ;
      LAYER met4 ;
        RECT 18.090000 198.790000 18.410000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 199.190000 18.410000 199.510000 ;
      LAYER met4 ;
        RECT 18.090000 199.190000 18.410000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090000 199.590000 18.410000 199.910000 ;
      LAYER met4 ;
        RECT 18.090000 199.590000 18.410000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 25.850000 18.695000 26.170000 ;
      LAYER met4 ;
        RECT 18.375000 25.850000 18.695000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 26.280000 18.695000 26.600000 ;
      LAYER met4 ;
        RECT 18.375000 26.280000 18.695000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 26.710000 18.695000 27.030000 ;
      LAYER met4 ;
        RECT 18.375000 26.710000 18.695000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 27.140000 18.695000 27.460000 ;
      LAYER met4 ;
        RECT 18.375000 27.140000 18.695000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 27.570000 18.695000 27.890000 ;
      LAYER met4 ;
        RECT 18.375000 27.570000 18.695000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 28.000000 18.695000 28.320000 ;
      LAYER met4 ;
        RECT 18.375000 28.000000 18.695000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 28.430000 18.695000 28.750000 ;
      LAYER met4 ;
        RECT 18.375000 28.430000 18.695000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 28.860000 18.695000 29.180000 ;
      LAYER met4 ;
        RECT 18.375000 28.860000 18.695000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 29.290000 18.695000 29.610000 ;
      LAYER met4 ;
        RECT 18.375000 29.290000 18.695000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 29.720000 18.695000 30.040000 ;
      LAYER met4 ;
        RECT 18.375000 29.720000 18.695000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 30.150000 18.695000 30.470000 ;
      LAYER met4 ;
        RECT 18.375000 30.150000 18.695000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 197.190000 18.815000 197.510000 ;
      LAYER met4 ;
        RECT 18.495000 197.190000 18.815000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 197.590000 18.815000 197.910000 ;
      LAYER met4 ;
        RECT 18.495000 197.590000 18.815000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 197.990000 18.815000 198.310000 ;
      LAYER met4 ;
        RECT 18.495000 197.990000 18.815000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 198.390000 18.815000 198.710000 ;
      LAYER met4 ;
        RECT 18.495000 198.390000 18.815000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 198.790000 18.815000 199.110000 ;
      LAYER met4 ;
        RECT 18.495000 198.790000 18.815000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 199.190000 18.815000 199.510000 ;
      LAYER met4 ;
        RECT 18.495000 199.190000 18.815000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 199.590000 18.815000 199.910000 ;
      LAYER met4 ;
        RECT 18.495000 199.590000 18.815000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 25.850000 19.100000 26.170000 ;
      LAYER met4 ;
        RECT 18.780000 25.850000 19.100000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 26.280000 19.100000 26.600000 ;
      LAYER met4 ;
        RECT 18.780000 26.280000 19.100000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 26.710000 19.100000 27.030000 ;
      LAYER met4 ;
        RECT 18.780000 26.710000 19.100000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 27.140000 19.100000 27.460000 ;
      LAYER met4 ;
        RECT 18.780000 27.140000 19.100000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 27.570000 19.100000 27.890000 ;
      LAYER met4 ;
        RECT 18.780000 27.570000 19.100000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 28.000000 19.100000 28.320000 ;
      LAYER met4 ;
        RECT 18.780000 28.000000 19.100000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 28.430000 19.100000 28.750000 ;
      LAYER met4 ;
        RECT 18.780000 28.430000 19.100000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 28.860000 19.100000 29.180000 ;
      LAYER met4 ;
        RECT 18.780000 28.860000 19.100000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 29.290000 19.100000 29.610000 ;
      LAYER met4 ;
        RECT 18.780000 29.290000 19.100000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 29.720000 19.100000 30.040000 ;
      LAYER met4 ;
        RECT 18.780000 29.720000 19.100000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 30.150000 19.100000 30.470000 ;
      LAYER met4 ;
        RECT 18.780000 30.150000 19.100000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 197.190000 19.220000 197.510000 ;
      LAYER met4 ;
        RECT 18.900000 197.190000 19.220000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 197.590000 19.220000 197.910000 ;
      LAYER met4 ;
        RECT 18.900000 197.590000 19.220000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 197.990000 19.220000 198.310000 ;
      LAYER met4 ;
        RECT 18.900000 197.990000 19.220000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 198.390000 19.220000 198.710000 ;
      LAYER met4 ;
        RECT 18.900000 198.390000 19.220000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 198.790000 19.220000 199.110000 ;
      LAYER met4 ;
        RECT 18.900000 198.790000 19.220000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 199.190000 19.220000 199.510000 ;
      LAYER met4 ;
        RECT 18.900000 199.190000 19.220000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900000 199.590000 19.220000 199.910000 ;
      LAYER met4 ;
        RECT 18.900000 199.590000 19.220000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 25.850000 19.505000 26.170000 ;
      LAYER met4 ;
        RECT 19.185000 25.850000 19.505000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 26.280000 19.505000 26.600000 ;
      LAYER met4 ;
        RECT 19.185000 26.280000 19.505000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 26.710000 19.505000 27.030000 ;
      LAYER met4 ;
        RECT 19.185000 26.710000 19.505000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 27.140000 19.505000 27.460000 ;
      LAYER met4 ;
        RECT 19.185000 27.140000 19.505000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 27.570000 19.505000 27.890000 ;
      LAYER met4 ;
        RECT 19.185000 27.570000 19.505000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 28.000000 19.505000 28.320000 ;
      LAYER met4 ;
        RECT 19.185000 28.000000 19.505000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 28.430000 19.505000 28.750000 ;
      LAYER met4 ;
        RECT 19.185000 28.430000 19.505000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 28.860000 19.505000 29.180000 ;
      LAYER met4 ;
        RECT 19.185000 28.860000 19.505000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 29.290000 19.505000 29.610000 ;
      LAYER met4 ;
        RECT 19.185000 29.290000 19.505000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 29.720000 19.505000 30.040000 ;
      LAYER met4 ;
        RECT 19.185000 29.720000 19.505000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 30.150000 19.505000 30.470000 ;
      LAYER met4 ;
        RECT 19.185000 30.150000 19.505000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 197.190000 19.625000 197.510000 ;
      LAYER met4 ;
        RECT 19.305000 197.190000 19.625000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 197.590000 19.625000 197.910000 ;
      LAYER met4 ;
        RECT 19.305000 197.590000 19.625000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 197.990000 19.625000 198.310000 ;
      LAYER met4 ;
        RECT 19.305000 197.990000 19.625000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 198.390000 19.625000 198.710000 ;
      LAYER met4 ;
        RECT 19.305000 198.390000 19.625000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 198.790000 19.625000 199.110000 ;
      LAYER met4 ;
        RECT 19.305000 198.790000 19.625000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 199.190000 19.625000 199.510000 ;
      LAYER met4 ;
        RECT 19.305000 199.190000 19.625000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305000 199.590000 19.625000 199.910000 ;
      LAYER met4 ;
        RECT 19.305000 199.590000 19.625000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 25.850000 19.910000 26.170000 ;
      LAYER met4 ;
        RECT 19.590000 25.850000 19.910000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 26.280000 19.910000 26.600000 ;
      LAYER met4 ;
        RECT 19.590000 26.280000 19.910000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 26.710000 19.910000 27.030000 ;
      LAYER met4 ;
        RECT 19.590000 26.710000 19.910000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 27.140000 19.910000 27.460000 ;
      LAYER met4 ;
        RECT 19.590000 27.140000 19.910000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 27.570000 19.910000 27.890000 ;
      LAYER met4 ;
        RECT 19.590000 27.570000 19.910000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 28.000000 19.910000 28.320000 ;
      LAYER met4 ;
        RECT 19.590000 28.000000 19.910000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 28.430000 19.910000 28.750000 ;
      LAYER met4 ;
        RECT 19.590000 28.430000 19.910000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 28.860000 19.910000 29.180000 ;
      LAYER met4 ;
        RECT 19.590000 28.860000 19.910000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 29.290000 19.910000 29.610000 ;
      LAYER met4 ;
        RECT 19.590000 29.290000 19.910000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 29.720000 19.910000 30.040000 ;
      LAYER met4 ;
        RECT 19.590000 29.720000 19.910000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 30.150000 19.910000 30.470000 ;
      LAYER met4 ;
        RECT 19.590000 30.150000 19.910000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 197.190000 20.030000 197.510000 ;
      LAYER met4 ;
        RECT 19.710000 197.190000 20.030000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 197.590000 20.030000 197.910000 ;
      LAYER met4 ;
        RECT 19.710000 197.590000 20.030000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 197.990000 20.030000 198.310000 ;
      LAYER met4 ;
        RECT 19.710000 197.990000 20.030000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 198.390000 20.030000 198.710000 ;
      LAYER met4 ;
        RECT 19.710000 198.390000 20.030000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 198.790000 20.030000 199.110000 ;
      LAYER met4 ;
        RECT 19.710000 198.790000 20.030000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 199.190000 20.030000 199.510000 ;
      LAYER met4 ;
        RECT 19.710000 199.190000 20.030000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710000 199.590000 20.030000 199.910000 ;
      LAYER met4 ;
        RECT 19.710000 199.590000 20.030000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 25.850000 20.315000 26.170000 ;
      LAYER met4 ;
        RECT 19.995000 25.850000 20.315000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 26.280000 20.315000 26.600000 ;
      LAYER met4 ;
        RECT 19.995000 26.280000 20.315000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 26.710000 20.315000 27.030000 ;
      LAYER met4 ;
        RECT 19.995000 26.710000 20.315000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 27.140000 20.315000 27.460000 ;
      LAYER met4 ;
        RECT 19.995000 27.140000 20.315000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 27.570000 20.315000 27.890000 ;
      LAYER met4 ;
        RECT 19.995000 27.570000 20.315000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 28.000000 20.315000 28.320000 ;
      LAYER met4 ;
        RECT 19.995000 28.000000 20.315000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 28.430000 20.315000 28.750000 ;
      LAYER met4 ;
        RECT 19.995000 28.430000 20.315000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 28.860000 20.315000 29.180000 ;
      LAYER met4 ;
        RECT 19.995000 28.860000 20.315000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 29.290000 20.315000 29.610000 ;
      LAYER met4 ;
        RECT 19.995000 29.290000 20.315000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 29.720000 20.315000 30.040000 ;
      LAYER met4 ;
        RECT 19.995000 29.720000 20.315000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 30.150000 20.315000 30.470000 ;
      LAYER met4 ;
        RECT 19.995000 30.150000 20.315000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 25.850000 2.485000 26.170000 ;
      LAYER met4 ;
        RECT 2.165000 25.850000 2.485000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 26.280000 2.485000 26.600000 ;
      LAYER met4 ;
        RECT 2.165000 26.280000 2.485000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 26.710000 2.485000 27.030000 ;
      LAYER met4 ;
        RECT 2.165000 26.710000 2.485000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 27.140000 2.485000 27.460000 ;
      LAYER met4 ;
        RECT 2.165000 27.140000 2.485000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 27.570000 2.485000 27.890000 ;
      LAYER met4 ;
        RECT 2.165000 27.570000 2.485000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 28.000000 2.485000 28.320000 ;
      LAYER met4 ;
        RECT 2.165000 28.000000 2.485000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 28.430000 2.485000 28.750000 ;
      LAYER met4 ;
        RECT 2.165000 28.430000 2.485000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 28.860000 2.485000 29.180000 ;
      LAYER met4 ;
        RECT 2.165000 28.860000 2.485000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 29.290000 2.485000 29.610000 ;
      LAYER met4 ;
        RECT 2.165000 29.290000 2.485000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 29.720000 2.485000 30.040000 ;
      LAYER met4 ;
        RECT 2.165000 29.720000 2.485000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 30.150000 2.485000 30.470000 ;
      LAYER met4 ;
        RECT 2.165000 30.150000 2.485000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 195.140000 2.545000 195.460000 ;
      LAYER met4 ;
        RECT 2.225000 195.140000 2.545000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 195.545000 2.545000 195.865000 ;
      LAYER met4 ;
        RECT 2.225000 195.545000 2.545000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 195.950000 2.545000 196.270000 ;
      LAYER met4 ;
        RECT 2.225000 195.950000 2.545000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 196.355000 2.545000 196.675000 ;
      LAYER met4 ;
        RECT 2.225000 196.355000 2.545000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 196.760000 2.545000 197.080000 ;
      LAYER met4 ;
        RECT 2.225000 196.760000 2.545000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 197.165000 2.545000 197.485000 ;
      LAYER met4 ;
        RECT 2.225000 197.165000 2.545000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 197.570000 2.545000 197.890000 ;
      LAYER met4 ;
        RECT 2.225000 197.570000 2.545000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 197.975000 2.545000 198.295000 ;
      LAYER met4 ;
        RECT 2.225000 197.975000 2.545000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 198.380000 2.545000 198.700000 ;
      LAYER met4 ;
        RECT 2.225000 198.380000 2.545000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 198.785000 2.545000 199.105000 ;
      LAYER met4 ;
        RECT 2.225000 198.785000 2.545000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 199.190000 2.545000 199.510000 ;
      LAYER met4 ;
        RECT 2.225000 199.190000 2.545000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225000 199.595000 2.545000 199.915000 ;
      LAYER met4 ;
        RECT 2.225000 199.595000 2.545000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 175.995000 2.485000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 176.395000 2.485000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 176.795000 2.485000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 177.195000 2.485000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 177.595000 2.485000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 177.995000 2.485000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 178.395000 2.485000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 178.795000 2.485000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 179.195000 2.485000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 179.595000 2.485000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 179.995000 2.485000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 180.395000 2.485000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 180.795000 2.485000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 181.195000 2.485000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 181.595000 2.485000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 181.995000 2.485000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 182.395000 2.485000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 182.795000 2.485000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 183.195000 2.485000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 183.595000 2.485000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 183.995000 2.485000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 184.395000 2.485000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 184.795000 2.485000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 185.195000 2.485000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 185.595000 2.485000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 185.995000 2.485000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 186.395000 2.485000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 186.795000 2.485000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 187.195000 2.485000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 187.595000 2.485000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 187.995000 2.485000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 188.395000 2.485000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 188.795000 2.485000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 189.195000 2.485000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 189.595000 2.485000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 189.995000 2.485000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 190.395000 2.485000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 190.795000 2.485000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 191.195000 2.485000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 191.595000 2.485000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 191.995000 2.485000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 192.395000 2.485000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 192.795000 2.485000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 193.195000 2.485000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 193.595000 2.485000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 193.995000 2.485000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 194.395000 2.485000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.285000 194.795000 2.485000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 25.850000 2.895000 26.170000 ;
      LAYER met4 ;
        RECT 2.575000 25.850000 2.895000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 26.280000 2.895000 26.600000 ;
      LAYER met4 ;
        RECT 2.575000 26.280000 2.895000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 26.710000 2.895000 27.030000 ;
      LAYER met4 ;
        RECT 2.575000 26.710000 2.895000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 27.140000 2.895000 27.460000 ;
      LAYER met4 ;
        RECT 2.575000 27.140000 2.895000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 27.570000 2.895000 27.890000 ;
      LAYER met4 ;
        RECT 2.575000 27.570000 2.895000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 28.000000 2.895000 28.320000 ;
      LAYER met4 ;
        RECT 2.575000 28.000000 2.895000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 28.430000 2.895000 28.750000 ;
      LAYER met4 ;
        RECT 2.575000 28.430000 2.895000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 28.860000 2.895000 29.180000 ;
      LAYER met4 ;
        RECT 2.575000 28.860000 2.895000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 29.290000 2.895000 29.610000 ;
      LAYER met4 ;
        RECT 2.575000 29.290000 2.895000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 29.720000 2.895000 30.040000 ;
      LAYER met4 ;
        RECT 2.575000 29.720000 2.895000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 30.150000 2.895000 30.470000 ;
      LAYER met4 ;
        RECT 2.575000 30.150000 2.895000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 195.140000 2.945000 195.460000 ;
      LAYER met4 ;
        RECT 2.625000 195.140000 2.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 195.545000 2.945000 195.865000 ;
      LAYER met4 ;
        RECT 2.625000 195.545000 2.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 195.950000 2.945000 196.270000 ;
      LAYER met4 ;
        RECT 2.625000 195.950000 2.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 196.355000 2.945000 196.675000 ;
      LAYER met4 ;
        RECT 2.625000 196.355000 2.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 196.760000 2.945000 197.080000 ;
      LAYER met4 ;
        RECT 2.625000 196.760000 2.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 197.165000 2.945000 197.485000 ;
      LAYER met4 ;
        RECT 2.625000 197.165000 2.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 197.570000 2.945000 197.890000 ;
      LAYER met4 ;
        RECT 2.625000 197.570000 2.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 197.975000 2.945000 198.295000 ;
      LAYER met4 ;
        RECT 2.625000 197.975000 2.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 198.380000 2.945000 198.700000 ;
      LAYER met4 ;
        RECT 2.625000 198.380000 2.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 198.785000 2.945000 199.105000 ;
      LAYER met4 ;
        RECT 2.625000 198.785000 2.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 199.190000 2.945000 199.510000 ;
      LAYER met4 ;
        RECT 2.625000 199.190000 2.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625000 199.595000 2.945000 199.915000 ;
      LAYER met4 ;
        RECT 2.625000 199.595000 2.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 175.995000 2.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 176.395000 2.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 176.795000 2.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 177.195000 2.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 177.595000 2.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 177.995000 2.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 178.395000 2.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 178.795000 2.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 179.195000 2.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 179.595000 2.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 179.995000 2.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 180.395000 2.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 180.795000 2.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 181.195000 2.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 181.595000 2.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 181.995000 2.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 182.395000 2.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 182.795000 2.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 183.195000 2.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 183.595000 2.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 183.995000 2.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 184.395000 2.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 184.795000 2.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 185.195000 2.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 185.595000 2.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 185.995000 2.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 186.395000 2.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 186.795000 2.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 187.195000 2.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 187.595000 2.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 187.995000 2.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 188.395000 2.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 188.795000 2.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 189.195000 2.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 189.595000 2.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 189.995000 2.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 190.395000 2.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 190.795000 2.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 191.195000 2.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 191.595000 2.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 191.995000 2.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 192.395000 2.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 192.795000 2.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 193.195000 2.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 193.595000 2.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 193.995000 2.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 194.395000 2.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.685000 194.795000 2.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 25.850000 3.305000 26.170000 ;
      LAYER met4 ;
        RECT 2.985000 25.850000 3.305000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 26.280000 3.305000 26.600000 ;
      LAYER met4 ;
        RECT 2.985000 26.280000 3.305000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 26.710000 3.305000 27.030000 ;
      LAYER met4 ;
        RECT 2.985000 26.710000 3.305000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 27.140000 3.305000 27.460000 ;
      LAYER met4 ;
        RECT 2.985000 27.140000 3.305000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 27.570000 3.305000 27.890000 ;
      LAYER met4 ;
        RECT 2.985000 27.570000 3.305000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 28.000000 3.305000 28.320000 ;
      LAYER met4 ;
        RECT 2.985000 28.000000 3.305000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 28.430000 3.305000 28.750000 ;
      LAYER met4 ;
        RECT 2.985000 28.430000 3.305000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 28.860000 3.305000 29.180000 ;
      LAYER met4 ;
        RECT 2.985000 28.860000 3.305000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 29.290000 3.305000 29.610000 ;
      LAYER met4 ;
        RECT 2.985000 29.290000 3.305000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 29.720000 3.305000 30.040000 ;
      LAYER met4 ;
        RECT 2.985000 29.720000 3.305000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 30.150000 3.305000 30.470000 ;
      LAYER met4 ;
        RECT 2.985000 30.150000 3.305000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 197.190000 20.435000 197.510000 ;
      LAYER met4 ;
        RECT 20.115000 197.190000 20.435000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 197.590000 20.435000 197.910000 ;
      LAYER met4 ;
        RECT 20.115000 197.590000 20.435000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 197.990000 20.435000 198.310000 ;
      LAYER met4 ;
        RECT 20.115000 197.990000 20.435000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 198.390000 20.435000 198.710000 ;
      LAYER met4 ;
        RECT 20.115000 198.390000 20.435000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 198.790000 20.435000 199.110000 ;
      LAYER met4 ;
        RECT 20.115000 198.790000 20.435000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 199.190000 20.435000 199.510000 ;
      LAYER met4 ;
        RECT 20.115000 199.190000 20.435000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115000 199.590000 20.435000 199.910000 ;
      LAYER met4 ;
        RECT 20.115000 199.590000 20.435000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 25.850000 20.720000 26.170000 ;
      LAYER met4 ;
        RECT 20.400000 25.850000 20.720000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 26.280000 20.720000 26.600000 ;
      LAYER met4 ;
        RECT 20.400000 26.280000 20.720000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 26.710000 20.720000 27.030000 ;
      LAYER met4 ;
        RECT 20.400000 26.710000 20.720000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 27.140000 20.720000 27.460000 ;
      LAYER met4 ;
        RECT 20.400000 27.140000 20.720000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 27.570000 20.720000 27.890000 ;
      LAYER met4 ;
        RECT 20.400000 27.570000 20.720000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 28.000000 20.720000 28.320000 ;
      LAYER met4 ;
        RECT 20.400000 28.000000 20.720000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 28.430000 20.720000 28.750000 ;
      LAYER met4 ;
        RECT 20.400000 28.430000 20.720000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 28.860000 20.720000 29.180000 ;
      LAYER met4 ;
        RECT 20.400000 28.860000 20.720000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 29.290000 20.720000 29.610000 ;
      LAYER met4 ;
        RECT 20.400000 29.290000 20.720000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 29.720000 20.720000 30.040000 ;
      LAYER met4 ;
        RECT 20.400000 29.720000 20.720000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 30.150000 20.720000 30.470000 ;
      LAYER met4 ;
        RECT 20.400000 30.150000 20.720000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 197.190000 20.840000 197.510000 ;
      LAYER met4 ;
        RECT 20.520000 197.190000 20.840000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 197.590000 20.840000 197.910000 ;
      LAYER met4 ;
        RECT 20.520000 197.590000 20.840000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 197.990000 20.840000 198.310000 ;
      LAYER met4 ;
        RECT 20.520000 197.990000 20.840000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 198.390000 20.840000 198.710000 ;
      LAYER met4 ;
        RECT 20.520000 198.390000 20.840000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 198.790000 20.840000 199.110000 ;
      LAYER met4 ;
        RECT 20.520000 198.790000 20.840000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 199.190000 20.840000 199.510000 ;
      LAYER met4 ;
        RECT 20.520000 199.190000 20.840000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520000 199.590000 20.840000 199.910000 ;
      LAYER met4 ;
        RECT 20.520000 199.590000 20.840000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 25.850000 21.125000 26.170000 ;
      LAYER met4 ;
        RECT 20.805000 25.850000 21.125000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 26.280000 21.125000 26.600000 ;
      LAYER met4 ;
        RECT 20.805000 26.280000 21.125000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 26.710000 21.125000 27.030000 ;
      LAYER met4 ;
        RECT 20.805000 26.710000 21.125000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 27.140000 21.125000 27.460000 ;
      LAYER met4 ;
        RECT 20.805000 27.140000 21.125000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 27.570000 21.125000 27.890000 ;
      LAYER met4 ;
        RECT 20.805000 27.570000 21.125000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 28.000000 21.125000 28.320000 ;
      LAYER met4 ;
        RECT 20.805000 28.000000 21.125000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 28.430000 21.125000 28.750000 ;
      LAYER met4 ;
        RECT 20.805000 28.430000 21.125000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 28.860000 21.125000 29.180000 ;
      LAYER met4 ;
        RECT 20.805000 28.860000 21.125000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 29.290000 21.125000 29.610000 ;
      LAYER met4 ;
        RECT 20.805000 29.290000 21.125000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 29.720000 21.125000 30.040000 ;
      LAYER met4 ;
        RECT 20.805000 29.720000 21.125000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 30.150000 21.125000 30.470000 ;
      LAYER met4 ;
        RECT 20.805000 30.150000 21.125000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 197.190000 21.245000 197.510000 ;
      LAYER met4 ;
        RECT 20.925000 197.190000 21.245000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 197.590000 21.245000 197.910000 ;
      LAYER met4 ;
        RECT 20.925000 197.590000 21.245000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 197.990000 21.245000 198.310000 ;
      LAYER met4 ;
        RECT 20.925000 197.990000 21.245000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 198.390000 21.245000 198.710000 ;
      LAYER met4 ;
        RECT 20.925000 198.390000 21.245000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 198.790000 21.245000 199.110000 ;
      LAYER met4 ;
        RECT 20.925000 198.790000 21.245000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 199.190000 21.245000 199.510000 ;
      LAYER met4 ;
        RECT 20.925000 199.190000 21.245000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925000 199.590000 21.245000 199.910000 ;
      LAYER met4 ;
        RECT 20.925000 199.590000 21.245000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 25.850000 21.530000 26.170000 ;
      LAYER met4 ;
        RECT 21.210000 25.850000 21.530000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 26.280000 21.530000 26.600000 ;
      LAYER met4 ;
        RECT 21.210000 26.280000 21.530000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 26.710000 21.530000 27.030000 ;
      LAYER met4 ;
        RECT 21.210000 26.710000 21.530000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 27.140000 21.530000 27.460000 ;
      LAYER met4 ;
        RECT 21.210000 27.140000 21.530000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 27.570000 21.530000 27.890000 ;
      LAYER met4 ;
        RECT 21.210000 27.570000 21.530000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 28.000000 21.530000 28.320000 ;
      LAYER met4 ;
        RECT 21.210000 28.000000 21.530000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 28.430000 21.530000 28.750000 ;
      LAYER met4 ;
        RECT 21.210000 28.430000 21.530000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 28.860000 21.530000 29.180000 ;
      LAYER met4 ;
        RECT 21.210000 28.860000 21.530000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 29.290000 21.530000 29.610000 ;
      LAYER met4 ;
        RECT 21.210000 29.290000 21.530000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 29.720000 21.530000 30.040000 ;
      LAYER met4 ;
        RECT 21.210000 29.720000 21.530000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 30.150000 21.530000 30.470000 ;
      LAYER met4 ;
        RECT 21.210000 30.150000 21.530000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 197.190000 21.650000 197.510000 ;
      LAYER met4 ;
        RECT 21.330000 197.190000 21.650000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 197.590000 21.650000 197.910000 ;
      LAYER met4 ;
        RECT 21.330000 197.590000 21.650000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 197.990000 21.650000 198.310000 ;
      LAYER met4 ;
        RECT 21.330000 197.990000 21.650000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 198.390000 21.650000 198.710000 ;
      LAYER met4 ;
        RECT 21.330000 198.390000 21.650000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 198.790000 21.650000 199.110000 ;
      LAYER met4 ;
        RECT 21.330000 198.790000 21.650000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 199.190000 21.650000 199.510000 ;
      LAYER met4 ;
        RECT 21.330000 199.190000 21.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330000 199.590000 21.650000 199.910000 ;
      LAYER met4 ;
        RECT 21.330000 199.590000 21.650000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 25.850000 21.935000 26.170000 ;
      LAYER met4 ;
        RECT 21.615000 25.850000 21.935000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 26.280000 21.935000 26.600000 ;
      LAYER met4 ;
        RECT 21.615000 26.280000 21.935000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 26.710000 21.935000 27.030000 ;
      LAYER met4 ;
        RECT 21.615000 26.710000 21.935000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 27.140000 21.935000 27.460000 ;
      LAYER met4 ;
        RECT 21.615000 27.140000 21.935000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 27.570000 21.935000 27.890000 ;
      LAYER met4 ;
        RECT 21.615000 27.570000 21.935000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 28.000000 21.935000 28.320000 ;
      LAYER met4 ;
        RECT 21.615000 28.000000 21.935000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 28.430000 21.935000 28.750000 ;
      LAYER met4 ;
        RECT 21.615000 28.430000 21.935000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 28.860000 21.935000 29.180000 ;
      LAYER met4 ;
        RECT 21.615000 28.860000 21.935000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 29.290000 21.935000 29.610000 ;
      LAYER met4 ;
        RECT 21.615000 29.290000 21.935000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 29.720000 21.935000 30.040000 ;
      LAYER met4 ;
        RECT 21.615000 29.720000 21.935000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 30.150000 21.935000 30.470000 ;
      LAYER met4 ;
        RECT 21.615000 30.150000 21.935000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 197.190000 22.055000 197.510000 ;
      LAYER met4 ;
        RECT 21.735000 197.190000 22.055000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 197.590000 22.055000 197.910000 ;
      LAYER met4 ;
        RECT 21.735000 197.590000 22.055000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 197.990000 22.055000 198.310000 ;
      LAYER met4 ;
        RECT 21.735000 197.990000 22.055000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 198.390000 22.055000 198.710000 ;
      LAYER met4 ;
        RECT 21.735000 198.390000 22.055000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 198.790000 22.055000 199.110000 ;
      LAYER met4 ;
        RECT 21.735000 198.790000 22.055000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 199.190000 22.055000 199.510000 ;
      LAYER met4 ;
        RECT 21.735000 199.190000 22.055000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735000 199.590000 22.055000 199.910000 ;
      LAYER met4 ;
        RECT 21.735000 199.590000 22.055000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 25.850000 22.340000 26.170000 ;
      LAYER met4 ;
        RECT 22.020000 25.850000 22.340000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 26.280000 22.340000 26.600000 ;
      LAYER met4 ;
        RECT 22.020000 26.280000 22.340000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 26.710000 22.340000 27.030000 ;
      LAYER met4 ;
        RECT 22.020000 26.710000 22.340000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 27.140000 22.340000 27.460000 ;
      LAYER met4 ;
        RECT 22.020000 27.140000 22.340000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 27.570000 22.340000 27.890000 ;
      LAYER met4 ;
        RECT 22.020000 27.570000 22.340000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 28.000000 22.340000 28.320000 ;
      LAYER met4 ;
        RECT 22.020000 28.000000 22.340000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 28.430000 22.340000 28.750000 ;
      LAYER met4 ;
        RECT 22.020000 28.430000 22.340000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 28.860000 22.340000 29.180000 ;
      LAYER met4 ;
        RECT 22.020000 28.860000 22.340000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 29.290000 22.340000 29.610000 ;
      LAYER met4 ;
        RECT 22.020000 29.290000 22.340000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 29.720000 22.340000 30.040000 ;
      LAYER met4 ;
        RECT 22.020000 29.720000 22.340000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 30.150000 22.340000 30.470000 ;
      LAYER met4 ;
        RECT 22.020000 30.150000 22.340000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 197.190000 22.460000 197.510000 ;
      LAYER met4 ;
        RECT 22.140000 197.190000 22.460000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 197.590000 22.460000 197.910000 ;
      LAYER met4 ;
        RECT 22.140000 197.590000 22.460000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 197.990000 22.460000 198.310000 ;
      LAYER met4 ;
        RECT 22.140000 197.990000 22.460000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 198.390000 22.460000 198.710000 ;
      LAYER met4 ;
        RECT 22.140000 198.390000 22.460000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 198.790000 22.460000 199.110000 ;
      LAYER met4 ;
        RECT 22.140000 198.790000 22.460000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 199.190000 22.460000 199.510000 ;
      LAYER met4 ;
        RECT 22.140000 199.190000 22.460000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140000 199.590000 22.460000 199.910000 ;
      LAYER met4 ;
        RECT 22.140000 199.590000 22.460000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 25.850000 22.745000 26.170000 ;
      LAYER met4 ;
        RECT 22.425000 25.850000 22.745000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 26.280000 22.745000 26.600000 ;
      LAYER met4 ;
        RECT 22.425000 26.280000 22.745000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 26.710000 22.745000 27.030000 ;
      LAYER met4 ;
        RECT 22.425000 26.710000 22.745000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 27.140000 22.745000 27.460000 ;
      LAYER met4 ;
        RECT 22.425000 27.140000 22.745000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 27.570000 22.745000 27.890000 ;
      LAYER met4 ;
        RECT 22.425000 27.570000 22.745000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 28.000000 22.745000 28.320000 ;
      LAYER met4 ;
        RECT 22.425000 28.000000 22.745000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 28.430000 22.745000 28.750000 ;
      LAYER met4 ;
        RECT 22.425000 28.430000 22.745000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 28.860000 22.745000 29.180000 ;
      LAYER met4 ;
        RECT 22.425000 28.860000 22.745000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 29.290000 22.745000 29.610000 ;
      LAYER met4 ;
        RECT 22.425000 29.290000 22.745000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 29.720000 22.745000 30.040000 ;
      LAYER met4 ;
        RECT 22.425000 29.720000 22.745000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 30.150000 22.745000 30.470000 ;
      LAYER met4 ;
        RECT 22.425000 30.150000 22.745000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 197.190000 22.865000 197.510000 ;
      LAYER met4 ;
        RECT 22.545000 197.190000 22.865000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 197.590000 22.865000 197.910000 ;
      LAYER met4 ;
        RECT 22.545000 197.590000 22.865000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 197.990000 22.865000 198.310000 ;
      LAYER met4 ;
        RECT 22.545000 197.990000 22.865000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 198.390000 22.865000 198.710000 ;
      LAYER met4 ;
        RECT 22.545000 198.390000 22.865000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 198.790000 22.865000 199.110000 ;
      LAYER met4 ;
        RECT 22.545000 198.790000 22.865000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 199.190000 22.865000 199.510000 ;
      LAYER met4 ;
        RECT 22.545000 199.190000 22.865000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 199.590000 22.865000 199.910000 ;
      LAYER met4 ;
        RECT 22.545000 199.590000 22.865000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 25.850000 23.150000 26.170000 ;
      LAYER met4 ;
        RECT 22.830000 25.850000 23.150000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 26.280000 23.150000 26.600000 ;
      LAYER met4 ;
        RECT 22.830000 26.280000 23.150000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 26.710000 23.150000 27.030000 ;
      LAYER met4 ;
        RECT 22.830000 26.710000 23.150000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 27.140000 23.150000 27.460000 ;
      LAYER met4 ;
        RECT 22.830000 27.140000 23.150000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 27.570000 23.150000 27.890000 ;
      LAYER met4 ;
        RECT 22.830000 27.570000 23.150000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 28.000000 23.150000 28.320000 ;
      LAYER met4 ;
        RECT 22.830000 28.000000 23.150000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 28.430000 23.150000 28.750000 ;
      LAYER met4 ;
        RECT 22.830000 28.430000 23.150000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 28.860000 23.150000 29.180000 ;
      LAYER met4 ;
        RECT 22.830000 28.860000 23.150000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 29.290000 23.150000 29.610000 ;
      LAYER met4 ;
        RECT 22.830000 29.290000 23.150000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 29.720000 23.150000 30.040000 ;
      LAYER met4 ;
        RECT 22.830000 29.720000 23.150000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 30.150000 23.150000 30.470000 ;
      LAYER met4 ;
        RECT 22.830000 30.150000 23.150000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 197.190000 23.270000 197.510000 ;
      LAYER met4 ;
        RECT 22.950000 197.190000 23.270000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 197.590000 23.270000 197.910000 ;
      LAYER met4 ;
        RECT 22.950000 197.590000 23.270000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 197.990000 23.270000 198.310000 ;
      LAYER met4 ;
        RECT 22.950000 197.990000 23.270000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 198.390000 23.270000 198.710000 ;
      LAYER met4 ;
        RECT 22.950000 198.390000 23.270000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 198.790000 23.270000 199.110000 ;
      LAYER met4 ;
        RECT 22.950000 198.790000 23.270000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 199.190000 23.270000 199.510000 ;
      LAYER met4 ;
        RECT 22.950000 199.190000 23.270000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 199.590000 23.270000 199.910000 ;
      LAYER met4 ;
        RECT 22.950000 199.590000 23.270000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 25.850000 23.555000 26.170000 ;
      LAYER met4 ;
        RECT 23.235000 25.850000 23.555000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 26.280000 23.555000 26.600000 ;
      LAYER met4 ;
        RECT 23.235000 26.280000 23.555000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 26.710000 23.555000 27.030000 ;
      LAYER met4 ;
        RECT 23.235000 26.710000 23.555000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 27.140000 23.555000 27.460000 ;
      LAYER met4 ;
        RECT 23.235000 27.140000 23.555000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 27.570000 23.555000 27.890000 ;
      LAYER met4 ;
        RECT 23.235000 27.570000 23.555000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 28.000000 23.555000 28.320000 ;
      LAYER met4 ;
        RECT 23.235000 28.000000 23.555000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 28.430000 23.555000 28.750000 ;
      LAYER met4 ;
        RECT 23.235000 28.430000 23.555000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 28.860000 23.555000 29.180000 ;
      LAYER met4 ;
        RECT 23.235000 28.860000 23.555000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 29.290000 23.555000 29.610000 ;
      LAYER met4 ;
        RECT 23.235000 29.290000 23.555000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 29.720000 23.555000 30.040000 ;
      LAYER met4 ;
        RECT 23.235000 29.720000 23.555000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 30.150000 23.555000 30.470000 ;
      LAYER met4 ;
        RECT 23.235000 30.150000 23.555000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 197.190000 23.675000 197.510000 ;
      LAYER met4 ;
        RECT 23.355000 197.190000 23.675000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 197.590000 23.675000 197.910000 ;
      LAYER met4 ;
        RECT 23.355000 197.590000 23.675000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 197.990000 23.675000 198.310000 ;
      LAYER met4 ;
        RECT 23.355000 197.990000 23.675000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 198.390000 23.675000 198.710000 ;
      LAYER met4 ;
        RECT 23.355000 198.390000 23.675000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 198.790000 23.675000 199.110000 ;
      LAYER met4 ;
        RECT 23.355000 198.790000 23.675000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 199.190000 23.675000 199.510000 ;
      LAYER met4 ;
        RECT 23.355000 199.190000 23.675000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355000 199.590000 23.675000 199.910000 ;
      LAYER met4 ;
        RECT 23.355000 199.590000 23.675000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 25.850000 23.960000 26.170000 ;
      LAYER met4 ;
        RECT 23.640000 25.850000 23.960000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 26.280000 23.960000 26.600000 ;
      LAYER met4 ;
        RECT 23.640000 26.280000 23.960000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 26.710000 23.960000 27.030000 ;
      LAYER met4 ;
        RECT 23.640000 26.710000 23.960000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 27.140000 23.960000 27.460000 ;
      LAYER met4 ;
        RECT 23.640000 27.140000 23.960000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 27.570000 23.960000 27.890000 ;
      LAYER met4 ;
        RECT 23.640000 27.570000 23.960000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 28.000000 23.960000 28.320000 ;
      LAYER met4 ;
        RECT 23.640000 28.000000 23.960000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 28.430000 23.960000 28.750000 ;
      LAYER met4 ;
        RECT 23.640000 28.430000 23.960000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 28.860000 23.960000 29.180000 ;
      LAYER met4 ;
        RECT 23.640000 28.860000 23.960000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 29.290000 23.960000 29.610000 ;
      LAYER met4 ;
        RECT 23.640000 29.290000 23.960000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 29.720000 23.960000 30.040000 ;
      LAYER met4 ;
        RECT 23.640000 29.720000 23.960000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 30.150000 23.960000 30.470000 ;
      LAYER met4 ;
        RECT 23.640000 30.150000 23.960000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 197.190000 24.080000 197.510000 ;
      LAYER met4 ;
        RECT 23.760000 197.190000 24.080000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 197.590000 24.080000 197.910000 ;
      LAYER met4 ;
        RECT 23.760000 197.590000 24.080000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 197.990000 24.080000 198.310000 ;
      LAYER met4 ;
        RECT 23.760000 197.990000 24.080000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 198.390000 24.080000 198.710000 ;
      LAYER met4 ;
        RECT 23.760000 198.390000 24.080000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 198.790000 24.080000 199.110000 ;
      LAYER met4 ;
        RECT 23.760000 198.790000 24.080000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 199.190000 24.080000 199.510000 ;
      LAYER met4 ;
        RECT 23.760000 199.190000 24.080000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760000 199.590000 24.080000 199.910000 ;
      LAYER met4 ;
        RECT 23.760000 199.590000 24.080000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 25.850000 24.365000 26.170000 ;
      LAYER met4 ;
        RECT 24.045000 25.850000 24.365000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 26.280000 24.365000 26.600000 ;
      LAYER met4 ;
        RECT 24.045000 26.280000 24.365000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 26.710000 24.365000 27.030000 ;
      LAYER met4 ;
        RECT 24.045000 26.710000 24.365000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 27.140000 24.365000 27.460000 ;
      LAYER met4 ;
        RECT 24.045000 27.140000 24.365000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 27.570000 24.365000 27.890000 ;
      LAYER met4 ;
        RECT 24.045000 27.570000 24.365000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 28.000000 24.365000 28.320000 ;
      LAYER met4 ;
        RECT 24.045000 28.000000 24.365000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 28.430000 24.365000 28.750000 ;
      LAYER met4 ;
        RECT 24.045000 28.430000 24.365000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 28.860000 24.365000 29.180000 ;
      LAYER met4 ;
        RECT 24.045000 28.860000 24.365000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 29.290000 24.365000 29.610000 ;
      LAYER met4 ;
        RECT 24.045000 29.290000 24.365000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 29.720000 24.365000 30.040000 ;
      LAYER met4 ;
        RECT 24.045000 29.720000 24.365000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 30.150000 24.365000 30.470000 ;
      LAYER met4 ;
        RECT 24.045000 30.150000 24.365000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 197.190000 24.485000 197.510000 ;
      LAYER met4 ;
        RECT 24.165000 197.190000 24.485000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 197.590000 24.485000 197.910000 ;
      LAYER met4 ;
        RECT 24.165000 197.590000 24.485000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 197.990000 24.485000 198.310000 ;
      LAYER met4 ;
        RECT 24.165000 197.990000 24.485000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 198.390000 24.485000 198.710000 ;
      LAYER met4 ;
        RECT 24.165000 198.390000 24.485000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 198.790000 24.485000 199.110000 ;
      LAYER met4 ;
        RECT 24.165000 198.790000 24.485000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 199.190000 24.485000 199.510000 ;
      LAYER met4 ;
        RECT 24.165000 199.190000 24.485000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165000 199.590000 24.485000 199.910000 ;
      LAYER met4 ;
        RECT 24.165000 199.590000 24.485000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 197.190000 24.890000 197.510000 ;
      LAYER met4 ;
        RECT 24.570000 197.190000 24.890000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 197.590000 24.890000 197.910000 ;
      LAYER met4 ;
        RECT 24.570000 197.590000 24.890000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 197.990000 24.890000 198.310000 ;
      LAYER met4 ;
        RECT 24.570000 197.990000 24.890000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 198.390000 24.890000 198.710000 ;
      LAYER met4 ;
        RECT 24.570000 198.390000 24.890000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 198.790000 24.890000 199.110000 ;
      LAYER met4 ;
        RECT 24.570000 198.790000 24.890000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 199.190000 24.890000 199.510000 ;
      LAYER met4 ;
        RECT 24.570000 199.190000 24.890000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570000 199.590000 24.890000 199.910000 ;
      LAYER met4 ;
        RECT 24.570000 199.590000 24.890000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 197.190000 25.295000 197.510000 ;
      LAYER met4 ;
        RECT 24.975000 197.190000 25.295000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 197.590000 25.295000 197.910000 ;
      LAYER met4 ;
        RECT 24.975000 197.590000 25.295000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 197.990000 25.295000 198.310000 ;
      LAYER met4 ;
        RECT 24.975000 197.990000 25.295000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 198.390000 25.295000 198.710000 ;
      LAYER met4 ;
        RECT 24.975000 198.390000 25.295000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 198.790000 25.295000 199.110000 ;
      LAYER met4 ;
        RECT 24.975000 198.790000 25.295000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 199.190000 25.295000 199.510000 ;
      LAYER met4 ;
        RECT 24.975000 199.190000 25.295000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975000 199.590000 25.295000 199.910000 ;
      LAYER met4 ;
        RECT 24.975000 199.590000 25.295000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 197.190000 25.700000 197.510000 ;
      LAYER met4 ;
        RECT 25.380000 197.190000 25.700000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 197.590000 25.700000 197.910000 ;
      LAYER met4 ;
        RECT 25.380000 197.590000 25.700000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 197.990000 25.700000 198.310000 ;
      LAYER met4 ;
        RECT 25.380000 197.990000 25.700000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 198.390000 25.700000 198.710000 ;
      LAYER met4 ;
        RECT 25.380000 198.390000 25.700000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 198.790000 25.700000 199.110000 ;
      LAYER met4 ;
        RECT 25.380000 198.790000 25.700000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 199.190000 25.700000 199.510000 ;
      LAYER met4 ;
        RECT 25.380000 199.190000 25.700000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380000 199.590000 25.700000 199.910000 ;
      LAYER met4 ;
        RECT 25.380000 199.590000 25.700000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 197.190000 26.105000 197.510000 ;
      LAYER met4 ;
        RECT 25.785000 197.190000 26.105000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 197.590000 26.105000 197.910000 ;
      LAYER met4 ;
        RECT 25.785000 197.590000 26.105000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 197.990000 26.105000 198.310000 ;
      LAYER met4 ;
        RECT 25.785000 197.990000 26.105000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 198.390000 26.105000 198.710000 ;
      LAYER met4 ;
        RECT 25.785000 198.390000 26.105000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 198.790000 26.105000 199.110000 ;
      LAYER met4 ;
        RECT 25.785000 198.790000 26.105000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 199.190000 26.105000 199.510000 ;
      LAYER met4 ;
        RECT 25.785000 199.190000 26.105000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785000 199.590000 26.105000 199.910000 ;
      LAYER met4 ;
        RECT 25.785000 199.590000 26.105000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 197.190000 26.510000 197.510000 ;
      LAYER met4 ;
        RECT 26.190000 197.190000 26.510000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 197.590000 26.510000 197.910000 ;
      LAYER met4 ;
        RECT 26.190000 197.590000 26.510000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 197.990000 26.510000 198.310000 ;
      LAYER met4 ;
        RECT 26.190000 197.990000 26.510000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 198.390000 26.510000 198.710000 ;
      LAYER met4 ;
        RECT 26.190000 198.390000 26.510000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 198.790000 26.510000 199.110000 ;
      LAYER met4 ;
        RECT 26.190000 198.790000 26.510000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 199.190000 26.510000 199.510000 ;
      LAYER met4 ;
        RECT 26.190000 199.190000 26.510000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190000 199.590000 26.510000 199.910000 ;
      LAYER met4 ;
        RECT 26.190000 199.590000 26.510000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 197.190000 26.915000 197.510000 ;
      LAYER met4 ;
        RECT 26.595000 197.190000 26.915000 197.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 197.590000 26.915000 197.910000 ;
      LAYER met4 ;
        RECT 26.595000 197.590000 26.915000 197.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 197.990000 26.915000 198.310000 ;
      LAYER met4 ;
        RECT 26.595000 197.990000 26.915000 198.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 198.390000 26.915000 198.710000 ;
      LAYER met4 ;
        RECT 26.595000 198.390000 26.915000 198.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 198.790000 26.915000 199.110000 ;
      LAYER met4 ;
        RECT 26.595000 198.790000 26.915000 199.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 199.190000 26.915000 199.510000 ;
      LAYER met4 ;
        RECT 26.595000 199.190000 26.915000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595000 199.590000 26.915000 199.910000 ;
      LAYER met4 ;
        RECT 26.595000 199.590000 26.915000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.000000 197.190000 37.060000 199.910000 ;
      LAYER met4 ;
        RECT 27.000000 197.190000 37.060000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 197.250000 27.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 197.650000 27.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 198.050000 27.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 198.450000 27.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 198.850000 27.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 199.250000 27.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.060000 199.650000 27.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 197.250000 27.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 197.650000 27.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 198.050000 27.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 198.450000 27.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 198.850000 27.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 199.250000 27.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.460000 199.650000 27.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 197.250000 28.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 197.650000 28.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 198.050000 28.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 198.450000 28.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 198.850000 28.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 199.250000 28.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.860000 199.650000 28.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 197.250000 28.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 197.650000 28.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 198.050000 28.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 198.450000 28.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 198.850000 28.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 199.250000 28.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.260000 199.650000 28.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 197.250000 28.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 197.650000 28.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 198.050000 28.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 198.450000 28.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 198.850000 28.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 199.250000 28.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.660000 199.650000 28.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 197.250000 29.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 197.650000 29.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 198.050000 29.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 198.450000 29.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 198.850000 29.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 199.250000 29.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.060000 199.650000 29.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 197.250000 29.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 197.650000 29.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 198.050000 29.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 198.450000 29.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 198.850000 29.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 199.250000 29.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.460000 199.650000 29.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 197.250000 30.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 197.650000 30.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 198.050000 30.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 198.450000 30.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 198.850000 30.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 199.250000 30.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.860000 199.650000 30.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 195.140000 3.345000 195.460000 ;
      LAYER met4 ;
        RECT 3.025000 195.140000 3.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 195.545000 3.345000 195.865000 ;
      LAYER met4 ;
        RECT 3.025000 195.545000 3.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 195.950000 3.345000 196.270000 ;
      LAYER met4 ;
        RECT 3.025000 195.950000 3.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 196.355000 3.345000 196.675000 ;
      LAYER met4 ;
        RECT 3.025000 196.355000 3.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 196.760000 3.345000 197.080000 ;
      LAYER met4 ;
        RECT 3.025000 196.760000 3.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 197.165000 3.345000 197.485000 ;
      LAYER met4 ;
        RECT 3.025000 197.165000 3.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 197.570000 3.345000 197.890000 ;
      LAYER met4 ;
        RECT 3.025000 197.570000 3.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 197.975000 3.345000 198.295000 ;
      LAYER met4 ;
        RECT 3.025000 197.975000 3.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 198.380000 3.345000 198.700000 ;
      LAYER met4 ;
        RECT 3.025000 198.380000 3.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 198.785000 3.345000 199.105000 ;
      LAYER met4 ;
        RECT 3.025000 198.785000 3.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 199.190000 3.345000 199.510000 ;
      LAYER met4 ;
        RECT 3.025000 199.190000 3.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 199.595000 3.345000 199.915000 ;
      LAYER met4 ;
        RECT 3.025000 199.595000 3.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 175.995000 3.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 176.395000 3.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 176.795000 3.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 177.195000 3.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 177.595000 3.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 177.995000 3.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 178.395000 3.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 178.795000 3.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 179.195000 3.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 179.595000 3.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 179.995000 3.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 180.395000 3.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 180.795000 3.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 181.195000 3.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 181.595000 3.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 181.995000 3.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 182.395000 3.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 182.795000 3.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 183.195000 3.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 183.595000 3.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 183.995000 3.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 184.395000 3.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 184.795000 3.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 185.195000 3.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 185.595000 3.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 185.995000 3.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 186.395000 3.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 186.795000 3.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 187.195000 3.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 187.595000 3.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 187.995000 3.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 188.395000 3.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 188.795000 3.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 189.195000 3.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 189.595000 3.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 189.995000 3.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 190.395000 3.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 190.795000 3.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 191.195000 3.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 191.595000 3.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 191.995000 3.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 192.395000 3.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 192.795000 3.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 193.195000 3.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 193.595000 3.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 193.995000 3.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 194.395000 3.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085000 194.795000 3.285000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 25.850000 3.710000 26.170000 ;
      LAYER met4 ;
        RECT 3.390000 25.850000 3.710000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 26.280000 3.710000 26.600000 ;
      LAYER met4 ;
        RECT 3.390000 26.280000 3.710000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 26.710000 3.710000 27.030000 ;
      LAYER met4 ;
        RECT 3.390000 26.710000 3.710000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 27.140000 3.710000 27.460000 ;
      LAYER met4 ;
        RECT 3.390000 27.140000 3.710000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 27.570000 3.710000 27.890000 ;
      LAYER met4 ;
        RECT 3.390000 27.570000 3.710000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 28.000000 3.710000 28.320000 ;
      LAYER met4 ;
        RECT 3.390000 28.000000 3.710000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 28.430000 3.710000 28.750000 ;
      LAYER met4 ;
        RECT 3.390000 28.430000 3.710000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 28.860000 3.710000 29.180000 ;
      LAYER met4 ;
        RECT 3.390000 28.860000 3.710000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 29.290000 3.710000 29.610000 ;
      LAYER met4 ;
        RECT 3.390000 29.290000 3.710000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 29.720000 3.710000 30.040000 ;
      LAYER met4 ;
        RECT 3.390000 29.720000 3.710000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 30.150000 3.710000 30.470000 ;
      LAYER met4 ;
        RECT 3.390000 30.150000 3.710000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 195.140000 3.745000 195.460000 ;
      LAYER met4 ;
        RECT 3.425000 195.140000 3.745000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 195.545000 3.745000 195.865000 ;
      LAYER met4 ;
        RECT 3.425000 195.545000 3.745000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 195.950000 3.745000 196.270000 ;
      LAYER met4 ;
        RECT 3.425000 195.950000 3.745000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 196.355000 3.745000 196.675000 ;
      LAYER met4 ;
        RECT 3.425000 196.355000 3.745000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 196.760000 3.745000 197.080000 ;
      LAYER met4 ;
        RECT 3.425000 196.760000 3.745000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 197.165000 3.745000 197.485000 ;
      LAYER met4 ;
        RECT 3.425000 197.165000 3.745000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 197.570000 3.745000 197.890000 ;
      LAYER met4 ;
        RECT 3.425000 197.570000 3.745000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 197.975000 3.745000 198.295000 ;
      LAYER met4 ;
        RECT 3.425000 197.975000 3.745000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 198.380000 3.745000 198.700000 ;
      LAYER met4 ;
        RECT 3.425000 198.380000 3.745000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 198.785000 3.745000 199.105000 ;
      LAYER met4 ;
        RECT 3.425000 198.785000 3.745000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 199.190000 3.745000 199.510000 ;
      LAYER met4 ;
        RECT 3.425000 199.190000 3.745000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425000 199.595000 3.745000 199.915000 ;
      LAYER met4 ;
        RECT 3.425000 199.595000 3.745000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 175.995000 3.685000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 176.395000 3.685000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 176.795000 3.685000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 177.195000 3.685000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 177.595000 3.685000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 177.995000 3.685000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 178.395000 3.685000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 178.795000 3.685000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 179.195000 3.685000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 179.595000 3.685000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 179.995000 3.685000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 180.395000 3.685000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 180.795000 3.685000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 181.195000 3.685000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 181.595000 3.685000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 181.995000 3.685000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 182.395000 3.685000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 182.795000 3.685000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 183.195000 3.685000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 183.595000 3.685000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 183.995000 3.685000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 184.395000 3.685000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 184.795000 3.685000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 185.195000 3.685000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 185.595000 3.685000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 185.995000 3.685000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 186.395000 3.685000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 186.795000 3.685000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 187.195000 3.685000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 187.595000 3.685000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 187.995000 3.685000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 188.395000 3.685000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 188.795000 3.685000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 189.195000 3.685000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 189.595000 3.685000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 189.995000 3.685000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 190.395000 3.685000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 190.795000 3.685000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 191.195000 3.685000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 191.595000 3.685000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 191.995000 3.685000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 192.395000 3.685000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 192.795000 3.685000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 193.195000 3.685000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 193.595000 3.685000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 193.995000 3.685000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 194.395000 3.685000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.485000 194.795000 3.685000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 25.850000 4.115000 26.170000 ;
      LAYER met4 ;
        RECT 3.795000 25.850000 4.115000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 26.280000 4.115000 26.600000 ;
      LAYER met4 ;
        RECT 3.795000 26.280000 4.115000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 26.710000 4.115000 27.030000 ;
      LAYER met4 ;
        RECT 3.795000 26.710000 4.115000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 27.140000 4.115000 27.460000 ;
      LAYER met4 ;
        RECT 3.795000 27.140000 4.115000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 27.570000 4.115000 27.890000 ;
      LAYER met4 ;
        RECT 3.795000 27.570000 4.115000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 28.000000 4.115000 28.320000 ;
      LAYER met4 ;
        RECT 3.795000 28.000000 4.115000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 28.430000 4.115000 28.750000 ;
      LAYER met4 ;
        RECT 3.795000 28.430000 4.115000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 28.860000 4.115000 29.180000 ;
      LAYER met4 ;
        RECT 3.795000 28.860000 4.115000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 29.290000 4.115000 29.610000 ;
      LAYER met4 ;
        RECT 3.795000 29.290000 4.115000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 29.720000 4.115000 30.040000 ;
      LAYER met4 ;
        RECT 3.795000 29.720000 4.115000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 30.150000 4.115000 30.470000 ;
      LAYER met4 ;
        RECT 3.795000 30.150000 4.115000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 195.140000 4.145000 195.460000 ;
      LAYER met4 ;
        RECT 3.825000 195.140000 4.145000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 195.545000 4.145000 195.865000 ;
      LAYER met4 ;
        RECT 3.825000 195.545000 4.145000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 195.950000 4.145000 196.270000 ;
      LAYER met4 ;
        RECT 3.825000 195.950000 4.145000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 196.355000 4.145000 196.675000 ;
      LAYER met4 ;
        RECT 3.825000 196.355000 4.145000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 196.760000 4.145000 197.080000 ;
      LAYER met4 ;
        RECT 3.825000 196.760000 4.145000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 197.165000 4.145000 197.485000 ;
      LAYER met4 ;
        RECT 3.825000 197.165000 4.145000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 197.570000 4.145000 197.890000 ;
      LAYER met4 ;
        RECT 3.825000 197.570000 4.145000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 197.975000 4.145000 198.295000 ;
      LAYER met4 ;
        RECT 3.825000 197.975000 4.145000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 198.380000 4.145000 198.700000 ;
      LAYER met4 ;
        RECT 3.825000 198.380000 4.145000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 198.785000 4.145000 199.105000 ;
      LAYER met4 ;
        RECT 3.825000 198.785000 4.145000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 199.190000 4.145000 199.510000 ;
      LAYER met4 ;
        RECT 3.825000 199.190000 4.145000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825000 199.595000 4.145000 199.915000 ;
      LAYER met4 ;
        RECT 3.825000 199.595000 4.145000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 175.995000 4.085000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 176.395000 4.085000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 176.795000 4.085000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 177.195000 4.085000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 177.595000 4.085000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 177.995000 4.085000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 178.395000 4.085000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 178.795000 4.085000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 179.195000 4.085000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 179.595000 4.085000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 179.995000 4.085000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 180.395000 4.085000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 180.795000 4.085000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 181.195000 4.085000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 181.595000 4.085000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 181.995000 4.085000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 182.395000 4.085000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 182.795000 4.085000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 183.195000 4.085000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 183.595000 4.085000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 183.995000 4.085000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 184.395000 4.085000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 184.795000 4.085000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 185.195000 4.085000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 185.595000 4.085000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 185.995000 4.085000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 186.395000 4.085000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 186.795000 4.085000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 187.195000 4.085000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 187.595000 4.085000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 187.995000 4.085000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 188.395000 4.085000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 188.795000 4.085000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 189.195000 4.085000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 189.595000 4.085000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 189.995000 4.085000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 190.395000 4.085000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 190.795000 4.085000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 191.195000 4.085000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 191.595000 4.085000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 191.995000 4.085000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 192.395000 4.085000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 192.795000 4.085000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 193.195000 4.085000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 193.595000 4.085000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 193.995000 4.085000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 194.395000 4.085000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.885000 194.795000 4.085000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 197.250000 30.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 197.650000 30.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 198.050000 30.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 198.450000 30.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 198.850000 30.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 199.250000 30.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.260000 199.650000 30.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 197.250000 30.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 197.650000 30.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 198.050000 30.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 198.450000 30.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 198.850000 30.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 199.250000 30.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.660000 199.650000 30.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 197.250000 31.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 197.650000 31.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 198.050000 31.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 198.450000 31.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 198.850000 31.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 199.250000 31.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.060000 199.650000 31.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 197.250000 31.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 197.650000 31.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 198.050000 31.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 198.450000 31.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 198.850000 31.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 199.250000 31.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.460000 199.650000 31.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 197.250000 32.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 197.650000 32.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 198.050000 32.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 198.450000 32.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 198.850000 32.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 199.250000 32.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.860000 199.650000 32.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 197.250000 32.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 197.650000 32.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 198.050000 32.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 198.450000 32.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 198.850000 32.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 199.250000 32.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.260000 199.650000 32.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 197.250000 32.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 197.650000 32.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 198.050000 32.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 198.450000 32.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 198.850000 32.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 199.250000 32.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.660000 199.650000 32.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 197.250000 33.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 197.650000 33.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 198.050000 33.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 198.450000 33.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 198.850000 33.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 199.250000 33.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.060000 199.650000 33.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 197.250000 33.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 197.650000 33.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 198.050000 33.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 198.450000 33.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 198.850000 33.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 199.250000 33.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.460000 199.650000 33.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 197.250000 34.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 197.650000 34.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 198.050000 34.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 198.450000 34.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 198.850000 34.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 199.250000 34.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.860000 199.650000 34.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 197.250000 34.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 197.650000 34.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 198.050000 34.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 198.450000 34.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 198.850000 34.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 199.250000 34.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.260000 199.650000 34.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 197.250000 34.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 197.650000 34.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 198.050000 34.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 198.450000 34.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 198.850000 34.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 199.250000 34.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.660000 199.650000 34.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 197.250000 35.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 197.650000 35.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 198.050000 35.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 198.450000 35.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 198.850000 35.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 199.250000 35.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.060000 199.650000 35.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 197.250000 35.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 197.650000 35.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 198.050000 35.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 198.450000 35.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 198.850000 35.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 199.250000 35.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.460000 199.650000 35.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 197.250000 36.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 197.650000 36.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 198.050000 36.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 198.450000 36.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 198.850000 36.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 199.250000 36.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.860000 199.650000 36.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 197.250000 36.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 197.650000 36.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 198.050000 36.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 198.450000 36.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 198.850000 36.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 199.250000 36.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.260000 199.650000 36.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.660000 197.250000 36.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.660000 197.650000 36.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.660000 198.050000 36.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.660000 198.450000 36.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.660000 198.850000 36.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.660000 199.250000 36.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 197.250000 37.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 197.650000 37.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 198.050000 37.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 198.450000 37.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 198.850000 37.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 199.250000 37.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.060000 199.650000 37.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.085000 197.190000 61.320000 199.910000 ;
      LAYER met4 ;
        RECT 37.085000 197.190000 61.320000 199.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 197.250000 37.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 197.650000 37.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 198.050000 37.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 198.450000 37.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 198.850000 37.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 199.250000 37.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.460000 199.650000 37.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 197.250000 38.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 197.650000 38.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 198.050000 38.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 198.450000 38.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 198.850000 38.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 199.250000 38.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.860000 199.650000 38.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 197.250000 38.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 197.650000 38.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 198.050000 38.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 198.450000 38.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 198.850000 38.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 199.250000 38.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.260000 199.650000 38.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 197.250000 38.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 197.650000 38.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 198.050000 38.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 198.450000 38.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 198.850000 38.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 199.250000 38.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.660000 199.650000 38.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 197.250000 39.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 197.650000 39.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 198.050000 39.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 198.450000 39.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 198.850000 39.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 199.250000 39.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.060000 199.650000 39.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 197.250000 39.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 197.650000 39.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 198.050000 39.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 198.450000 39.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 198.850000 39.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 199.250000 39.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.460000 199.650000 39.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 197.250000 40.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 197.650000 40.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 198.050000 40.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 198.450000 40.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 198.850000 40.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 199.250000 40.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.860000 199.650000 40.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 25.850000 4.520000 26.170000 ;
      LAYER met4 ;
        RECT 4.200000 25.850000 4.520000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 26.280000 4.520000 26.600000 ;
      LAYER met4 ;
        RECT 4.200000 26.280000 4.520000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 26.710000 4.520000 27.030000 ;
      LAYER met4 ;
        RECT 4.200000 26.710000 4.520000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 27.140000 4.520000 27.460000 ;
      LAYER met4 ;
        RECT 4.200000 27.140000 4.520000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 27.570000 4.520000 27.890000 ;
      LAYER met4 ;
        RECT 4.200000 27.570000 4.520000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 28.000000 4.520000 28.320000 ;
      LAYER met4 ;
        RECT 4.200000 28.000000 4.520000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 28.430000 4.520000 28.750000 ;
      LAYER met4 ;
        RECT 4.200000 28.430000 4.520000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 28.860000 4.520000 29.180000 ;
      LAYER met4 ;
        RECT 4.200000 28.860000 4.520000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 29.290000 4.520000 29.610000 ;
      LAYER met4 ;
        RECT 4.200000 29.290000 4.520000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 29.720000 4.520000 30.040000 ;
      LAYER met4 ;
        RECT 4.200000 29.720000 4.520000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 30.150000 4.520000 30.470000 ;
      LAYER met4 ;
        RECT 4.200000 30.150000 4.520000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 195.140000 4.545000 195.460000 ;
      LAYER met4 ;
        RECT 4.225000 195.140000 4.545000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 195.545000 4.545000 195.865000 ;
      LAYER met4 ;
        RECT 4.225000 195.545000 4.545000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 195.950000 4.545000 196.270000 ;
      LAYER met4 ;
        RECT 4.225000 195.950000 4.545000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 196.355000 4.545000 196.675000 ;
      LAYER met4 ;
        RECT 4.225000 196.355000 4.545000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 196.760000 4.545000 197.080000 ;
      LAYER met4 ;
        RECT 4.225000 196.760000 4.545000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 197.165000 4.545000 197.485000 ;
      LAYER met4 ;
        RECT 4.225000 197.165000 4.545000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 197.570000 4.545000 197.890000 ;
      LAYER met4 ;
        RECT 4.225000 197.570000 4.545000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 197.975000 4.545000 198.295000 ;
      LAYER met4 ;
        RECT 4.225000 197.975000 4.545000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 198.380000 4.545000 198.700000 ;
      LAYER met4 ;
        RECT 4.225000 198.380000 4.545000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 198.785000 4.545000 199.105000 ;
      LAYER met4 ;
        RECT 4.225000 198.785000 4.545000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 199.190000 4.545000 199.510000 ;
      LAYER met4 ;
        RECT 4.225000 199.190000 4.545000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225000 199.595000 4.545000 199.915000 ;
      LAYER met4 ;
        RECT 4.225000 199.595000 4.545000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 175.995000 4.485000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 176.395000 4.485000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 176.795000 4.485000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 177.195000 4.485000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 177.595000 4.485000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 177.995000 4.485000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 178.395000 4.485000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 178.795000 4.485000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 179.195000 4.485000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 179.595000 4.485000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 179.995000 4.485000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 180.395000 4.485000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 180.795000 4.485000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 181.195000 4.485000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 181.595000 4.485000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 181.995000 4.485000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 182.395000 4.485000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 182.795000 4.485000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 183.195000 4.485000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 183.595000 4.485000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 183.995000 4.485000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 184.395000 4.485000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 184.795000 4.485000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 185.195000 4.485000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 185.595000 4.485000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 185.995000 4.485000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 186.395000 4.485000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 186.795000 4.485000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 187.195000 4.485000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 187.595000 4.485000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 187.995000 4.485000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 188.395000 4.485000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 188.795000 4.485000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 189.195000 4.485000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 189.595000 4.485000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 189.995000 4.485000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 190.395000 4.485000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 190.795000 4.485000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 191.195000 4.485000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 191.595000 4.485000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 191.995000 4.485000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 192.395000 4.485000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 192.795000 4.485000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 193.195000 4.485000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 193.595000 4.485000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 193.995000 4.485000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 194.395000 4.485000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.285000 194.795000 4.485000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 25.850000 4.925000 26.170000 ;
      LAYER met4 ;
        RECT 4.605000 25.850000 4.925000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 26.280000 4.925000 26.600000 ;
      LAYER met4 ;
        RECT 4.605000 26.280000 4.925000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 26.710000 4.925000 27.030000 ;
      LAYER met4 ;
        RECT 4.605000 26.710000 4.925000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 27.140000 4.925000 27.460000 ;
      LAYER met4 ;
        RECT 4.605000 27.140000 4.925000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 27.570000 4.925000 27.890000 ;
      LAYER met4 ;
        RECT 4.605000 27.570000 4.925000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 28.000000 4.925000 28.320000 ;
      LAYER met4 ;
        RECT 4.605000 28.000000 4.925000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 28.430000 4.925000 28.750000 ;
      LAYER met4 ;
        RECT 4.605000 28.430000 4.925000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 28.860000 4.925000 29.180000 ;
      LAYER met4 ;
        RECT 4.605000 28.860000 4.925000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 29.290000 4.925000 29.610000 ;
      LAYER met4 ;
        RECT 4.605000 29.290000 4.925000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 29.720000 4.925000 30.040000 ;
      LAYER met4 ;
        RECT 4.605000 29.720000 4.925000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 30.150000 4.925000 30.470000 ;
      LAYER met4 ;
        RECT 4.605000 30.150000 4.925000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 195.140000 4.945000 195.460000 ;
      LAYER met4 ;
        RECT 4.625000 195.140000 4.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 195.545000 4.945000 195.865000 ;
      LAYER met4 ;
        RECT 4.625000 195.545000 4.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 195.950000 4.945000 196.270000 ;
      LAYER met4 ;
        RECT 4.625000 195.950000 4.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 196.355000 4.945000 196.675000 ;
      LAYER met4 ;
        RECT 4.625000 196.355000 4.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 196.760000 4.945000 197.080000 ;
      LAYER met4 ;
        RECT 4.625000 196.760000 4.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 197.165000 4.945000 197.485000 ;
      LAYER met4 ;
        RECT 4.625000 197.165000 4.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 197.570000 4.945000 197.890000 ;
      LAYER met4 ;
        RECT 4.625000 197.570000 4.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 197.975000 4.945000 198.295000 ;
      LAYER met4 ;
        RECT 4.625000 197.975000 4.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 198.380000 4.945000 198.700000 ;
      LAYER met4 ;
        RECT 4.625000 198.380000 4.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 198.785000 4.945000 199.105000 ;
      LAYER met4 ;
        RECT 4.625000 198.785000 4.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 199.190000 4.945000 199.510000 ;
      LAYER met4 ;
        RECT 4.625000 199.190000 4.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625000 199.595000 4.945000 199.915000 ;
      LAYER met4 ;
        RECT 4.625000 199.595000 4.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 175.995000 4.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 176.395000 4.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 176.795000 4.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 177.195000 4.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 177.595000 4.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 177.995000 4.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 178.395000 4.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 178.795000 4.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 179.195000 4.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 179.595000 4.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 179.995000 4.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 180.395000 4.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 180.795000 4.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 181.195000 4.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 181.595000 4.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 181.995000 4.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 182.395000 4.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 182.795000 4.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 183.195000 4.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 183.595000 4.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 183.995000 4.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 184.395000 4.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 184.795000 4.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 185.195000 4.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 185.595000 4.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 185.995000 4.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 186.395000 4.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 186.795000 4.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 187.195000 4.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 187.595000 4.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 187.995000 4.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 188.395000 4.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 188.795000 4.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 189.195000 4.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 189.595000 4.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 189.995000 4.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 190.395000 4.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 190.795000 4.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 191.195000 4.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 191.595000 4.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 191.995000 4.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 192.395000 4.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 192.795000 4.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 193.195000 4.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 193.595000 4.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 193.995000 4.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 194.395000 4.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.685000 194.795000 4.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 197.250000 40.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 197.650000 40.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 198.050000 40.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 198.450000 40.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 198.850000 40.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 199.250000 40.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.260000 199.650000 40.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 197.250000 40.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 197.650000 40.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 198.050000 40.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 198.450000 40.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 198.850000 40.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 199.250000 40.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.660000 199.650000 40.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 197.250000 41.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 197.650000 41.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 198.050000 41.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 198.450000 41.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 198.850000 41.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 199.250000 41.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.060000 199.650000 41.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 197.250000 41.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 197.650000 41.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 198.050000 41.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 198.450000 41.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 198.850000 41.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 199.250000 41.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.460000 199.650000 41.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 197.250000 42.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 197.650000 42.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 198.050000 42.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 198.450000 42.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 198.850000 42.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 199.250000 42.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.860000 199.650000 42.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 197.250000 42.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 197.650000 42.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 198.050000 42.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 198.450000 42.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 198.850000 42.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 199.250000 42.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.260000 199.650000 42.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 197.250000 42.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 197.650000 42.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 198.050000 42.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 198.450000 42.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 198.850000 42.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 199.250000 42.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.660000 199.650000 42.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 197.250000 43.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 197.650000 43.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 198.050000 43.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 198.450000 43.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 198.850000 43.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 199.250000 43.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.060000 199.650000 43.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 197.250000 43.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 197.650000 43.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 198.050000 43.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 198.450000 43.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 198.850000 43.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 199.250000 43.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.460000 199.650000 43.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 197.250000 44.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 197.650000 44.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 198.050000 44.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 198.450000 44.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 198.850000 44.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 199.250000 44.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.860000 199.650000 44.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 197.250000 44.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 197.650000 44.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 198.050000 44.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 198.450000 44.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 198.850000 44.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 199.250000 44.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.260000 199.650000 44.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 197.250000 44.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 197.650000 44.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 198.050000 44.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 198.450000 44.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 198.850000 44.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 199.250000 44.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.660000 199.650000 44.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 197.250000 45.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 197.650000 45.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 198.050000 45.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 198.450000 45.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 198.850000 45.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 199.250000 45.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 199.650000 45.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 197.250000 45.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 197.650000 45.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 198.050000 45.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 198.450000 45.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 198.850000 45.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 199.250000 45.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.460000 199.650000 45.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 197.250000 46.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 197.650000 46.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 198.050000 46.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 198.450000 46.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 198.850000 46.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 199.250000 46.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 199.650000 46.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 197.250000 46.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 197.650000 46.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 198.050000 46.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 198.450000 46.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 198.850000 46.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 199.250000 46.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.260000 199.650000 46.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 197.250000 46.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 197.650000 46.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 198.050000 46.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 198.450000 46.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 198.850000 46.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 199.250000 46.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.660000 199.650000 46.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 197.250000 47.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 197.650000 47.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 198.050000 47.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 198.450000 47.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 198.850000 47.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 199.250000 47.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 199.650000 47.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 197.250000 47.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 197.650000 47.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 198.050000 47.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 198.450000 47.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 198.850000 47.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 199.250000 47.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.460000 199.650000 47.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 197.250000 48.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 197.650000 48.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 198.050000 48.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 198.450000 48.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 198.850000 48.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 199.250000 48.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.860000 199.650000 48.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 197.250000 48.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 197.650000 48.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 198.050000 48.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 198.450000 48.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 198.850000 48.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 199.250000 48.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 199.650000 48.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 197.250000 48.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 197.650000 48.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 198.050000 48.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 198.450000 48.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 198.850000 48.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 199.250000 48.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.660000 199.650000 48.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 197.250000 49.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 197.650000 49.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 198.050000 49.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 198.450000 49.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 198.850000 49.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 199.250000 49.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.060000 199.650000 49.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 197.250000 49.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 197.650000 49.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 198.050000 49.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 198.450000 49.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 198.850000 49.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 199.250000 49.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 199.650000 49.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 197.250000 50.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 197.650000 50.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 198.050000 50.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 198.450000 50.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 198.850000 50.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 199.250000 50.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.860000 199.650000 50.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 25.850000 5.330000 26.170000 ;
      LAYER met4 ;
        RECT 5.010000 25.850000 5.330000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 26.280000 5.330000 26.600000 ;
      LAYER met4 ;
        RECT 5.010000 26.280000 5.330000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 26.710000 5.330000 27.030000 ;
      LAYER met4 ;
        RECT 5.010000 26.710000 5.330000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 27.140000 5.330000 27.460000 ;
      LAYER met4 ;
        RECT 5.010000 27.140000 5.330000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 27.570000 5.330000 27.890000 ;
      LAYER met4 ;
        RECT 5.010000 27.570000 5.330000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 28.000000 5.330000 28.320000 ;
      LAYER met4 ;
        RECT 5.010000 28.000000 5.330000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 28.430000 5.330000 28.750000 ;
      LAYER met4 ;
        RECT 5.010000 28.430000 5.330000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 28.860000 5.330000 29.180000 ;
      LAYER met4 ;
        RECT 5.010000 28.860000 5.330000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 29.290000 5.330000 29.610000 ;
      LAYER met4 ;
        RECT 5.010000 29.290000 5.330000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 29.720000 5.330000 30.040000 ;
      LAYER met4 ;
        RECT 5.010000 29.720000 5.330000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 30.150000 5.330000 30.470000 ;
      LAYER met4 ;
        RECT 5.010000 30.150000 5.330000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 195.140000 5.345000 195.460000 ;
      LAYER met4 ;
        RECT 5.025000 195.140000 5.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 195.545000 5.345000 195.865000 ;
      LAYER met4 ;
        RECT 5.025000 195.545000 5.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 195.950000 5.345000 196.270000 ;
      LAYER met4 ;
        RECT 5.025000 195.950000 5.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 196.355000 5.345000 196.675000 ;
      LAYER met4 ;
        RECT 5.025000 196.355000 5.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 196.760000 5.345000 197.080000 ;
      LAYER met4 ;
        RECT 5.025000 196.760000 5.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 197.165000 5.345000 197.485000 ;
      LAYER met4 ;
        RECT 5.025000 197.165000 5.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 197.570000 5.345000 197.890000 ;
      LAYER met4 ;
        RECT 5.025000 197.570000 5.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 197.975000 5.345000 198.295000 ;
      LAYER met4 ;
        RECT 5.025000 197.975000 5.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 198.380000 5.345000 198.700000 ;
      LAYER met4 ;
        RECT 5.025000 198.380000 5.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 198.785000 5.345000 199.105000 ;
      LAYER met4 ;
        RECT 5.025000 198.785000 5.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 199.190000 5.345000 199.510000 ;
      LAYER met4 ;
        RECT 5.025000 199.190000 5.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025000 199.595000 5.345000 199.915000 ;
      LAYER met4 ;
        RECT 5.025000 199.595000 5.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 175.995000 5.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 176.395000 5.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 176.795000 5.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 177.195000 5.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 177.595000 5.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 177.995000 5.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 178.395000 5.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 178.795000 5.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 179.195000 5.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 179.595000 5.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 179.995000 5.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 180.395000 5.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 180.795000 5.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 181.195000 5.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 181.595000 5.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 181.995000 5.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 182.395000 5.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 182.795000 5.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 183.195000 5.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 183.595000 5.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 183.995000 5.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 184.395000 5.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 184.795000 5.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 185.195000 5.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 185.595000 5.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 185.995000 5.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 186.395000 5.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 186.795000 5.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 187.195000 5.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 187.595000 5.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 187.995000 5.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 188.395000 5.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 188.795000 5.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 189.195000 5.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 189.595000 5.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 189.995000 5.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 190.395000 5.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 190.795000 5.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 191.195000 5.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 191.595000 5.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 191.995000 5.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 192.395000 5.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 192.795000 5.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 193.195000 5.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 193.595000 5.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 193.995000 5.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 194.395000 5.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 194.795000 5.285000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 25.850000 5.735000 26.170000 ;
      LAYER met4 ;
        RECT 5.415000 25.850000 5.735000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 26.280000 5.735000 26.600000 ;
      LAYER met4 ;
        RECT 5.415000 26.280000 5.735000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 26.710000 5.735000 27.030000 ;
      LAYER met4 ;
        RECT 5.415000 26.710000 5.735000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 27.140000 5.735000 27.460000 ;
      LAYER met4 ;
        RECT 5.415000 27.140000 5.735000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 27.570000 5.735000 27.890000 ;
      LAYER met4 ;
        RECT 5.415000 27.570000 5.735000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 28.000000 5.735000 28.320000 ;
      LAYER met4 ;
        RECT 5.415000 28.000000 5.735000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 28.430000 5.735000 28.750000 ;
      LAYER met4 ;
        RECT 5.415000 28.430000 5.735000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 28.860000 5.735000 29.180000 ;
      LAYER met4 ;
        RECT 5.415000 28.860000 5.735000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 29.290000 5.735000 29.610000 ;
      LAYER met4 ;
        RECT 5.415000 29.290000 5.735000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 29.720000 5.735000 30.040000 ;
      LAYER met4 ;
        RECT 5.415000 29.720000 5.735000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 30.150000 5.735000 30.470000 ;
      LAYER met4 ;
        RECT 5.415000 30.150000 5.735000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 195.140000 5.745000 195.460000 ;
      LAYER met4 ;
        RECT 5.425000 195.140000 5.745000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 195.545000 5.745000 195.865000 ;
      LAYER met4 ;
        RECT 5.425000 195.545000 5.745000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 195.950000 5.745000 196.270000 ;
      LAYER met4 ;
        RECT 5.425000 195.950000 5.745000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 196.355000 5.745000 196.675000 ;
      LAYER met4 ;
        RECT 5.425000 196.355000 5.745000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 196.760000 5.745000 197.080000 ;
      LAYER met4 ;
        RECT 5.425000 196.760000 5.745000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 197.165000 5.745000 197.485000 ;
      LAYER met4 ;
        RECT 5.425000 197.165000 5.745000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 197.570000 5.745000 197.890000 ;
      LAYER met4 ;
        RECT 5.425000 197.570000 5.745000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 197.975000 5.745000 198.295000 ;
      LAYER met4 ;
        RECT 5.425000 197.975000 5.745000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 198.380000 5.745000 198.700000 ;
      LAYER met4 ;
        RECT 5.425000 198.380000 5.745000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 198.785000 5.745000 199.105000 ;
      LAYER met4 ;
        RECT 5.425000 198.785000 5.745000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 199.190000 5.745000 199.510000 ;
      LAYER met4 ;
        RECT 5.425000 199.190000 5.745000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425000 199.595000 5.745000 199.915000 ;
      LAYER met4 ;
        RECT 5.425000 199.595000 5.745000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 175.995000 5.685000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 176.395000 5.685000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 176.795000 5.685000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 177.195000 5.685000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 177.595000 5.685000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 177.995000 5.685000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 178.395000 5.685000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 178.795000 5.685000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 179.195000 5.685000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 179.595000 5.685000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 179.995000 5.685000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 180.395000 5.685000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 180.795000 5.685000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 181.195000 5.685000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 181.595000 5.685000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 181.995000 5.685000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 182.395000 5.685000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 182.795000 5.685000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 183.195000 5.685000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 183.595000 5.685000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 183.995000 5.685000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 184.395000 5.685000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 184.795000 5.685000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 185.195000 5.685000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 185.595000 5.685000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 185.995000 5.685000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 186.395000 5.685000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 186.795000 5.685000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 187.195000 5.685000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 187.595000 5.685000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 187.995000 5.685000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 188.395000 5.685000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 188.795000 5.685000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 189.195000 5.685000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 189.595000 5.685000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 189.995000 5.685000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 190.395000 5.685000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 190.795000 5.685000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 191.195000 5.685000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 191.595000 5.685000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 191.995000 5.685000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 192.395000 5.685000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 192.795000 5.685000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 193.195000 5.685000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 193.595000 5.685000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 193.995000 5.685000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 194.395000 5.685000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.485000 194.795000 5.685000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 25.850000 6.140000 26.170000 ;
      LAYER met4 ;
        RECT 5.820000 25.850000 6.140000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 26.280000 6.140000 26.600000 ;
      LAYER met4 ;
        RECT 5.820000 26.280000 6.140000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 26.710000 6.140000 27.030000 ;
      LAYER met4 ;
        RECT 5.820000 26.710000 6.140000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 27.140000 6.140000 27.460000 ;
      LAYER met4 ;
        RECT 5.820000 27.140000 6.140000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 27.570000 6.140000 27.890000 ;
      LAYER met4 ;
        RECT 5.820000 27.570000 6.140000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 28.000000 6.140000 28.320000 ;
      LAYER met4 ;
        RECT 5.820000 28.000000 6.140000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 28.430000 6.140000 28.750000 ;
      LAYER met4 ;
        RECT 5.820000 28.430000 6.140000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 28.860000 6.140000 29.180000 ;
      LAYER met4 ;
        RECT 5.820000 28.860000 6.140000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 29.290000 6.140000 29.610000 ;
      LAYER met4 ;
        RECT 5.820000 29.290000 6.140000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 29.720000 6.140000 30.040000 ;
      LAYER met4 ;
        RECT 5.820000 29.720000 6.140000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 30.150000 6.140000 30.470000 ;
      LAYER met4 ;
        RECT 5.820000 30.150000 6.140000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 195.140000 6.145000 195.460000 ;
      LAYER met4 ;
        RECT 5.825000 195.140000 6.145000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 195.545000 6.145000 195.865000 ;
      LAYER met4 ;
        RECT 5.825000 195.545000 6.145000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 195.950000 6.145000 196.270000 ;
      LAYER met4 ;
        RECT 5.825000 195.950000 6.145000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 196.355000 6.145000 196.675000 ;
      LAYER met4 ;
        RECT 5.825000 196.355000 6.145000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 196.760000 6.145000 197.080000 ;
      LAYER met4 ;
        RECT 5.825000 196.760000 6.145000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 197.165000 6.145000 197.485000 ;
      LAYER met4 ;
        RECT 5.825000 197.165000 6.145000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 197.570000 6.145000 197.890000 ;
      LAYER met4 ;
        RECT 5.825000 197.570000 6.145000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 197.975000 6.145000 198.295000 ;
      LAYER met4 ;
        RECT 5.825000 197.975000 6.145000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 198.380000 6.145000 198.700000 ;
      LAYER met4 ;
        RECT 5.825000 198.380000 6.145000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 198.785000 6.145000 199.105000 ;
      LAYER met4 ;
        RECT 5.825000 198.785000 6.145000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 199.190000 6.145000 199.510000 ;
      LAYER met4 ;
        RECT 5.825000 199.190000 6.145000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 199.595000 6.145000 199.915000 ;
      LAYER met4 ;
        RECT 5.825000 199.595000 6.145000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 175.995000 6.085000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 176.395000 6.085000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 176.795000 6.085000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 177.195000 6.085000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 177.595000 6.085000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 177.995000 6.085000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 178.395000 6.085000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 178.795000 6.085000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 179.195000 6.085000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 179.595000 6.085000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 179.995000 6.085000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 180.395000 6.085000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 180.795000 6.085000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 181.195000 6.085000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 181.595000 6.085000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 181.995000 6.085000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 182.395000 6.085000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 182.795000 6.085000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 183.195000 6.085000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 183.595000 6.085000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 183.995000 6.085000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 184.395000 6.085000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 184.795000 6.085000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 185.195000 6.085000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 185.595000 6.085000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 185.995000 6.085000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 186.395000 6.085000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 186.795000 6.085000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 187.195000 6.085000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 187.595000 6.085000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 187.995000 6.085000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 188.395000 6.085000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 188.795000 6.085000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 189.195000 6.085000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 189.595000 6.085000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 189.995000 6.085000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 190.395000 6.085000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 190.795000 6.085000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 191.195000 6.085000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 191.595000 6.085000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 191.995000 6.085000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 192.395000 6.085000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 192.795000 6.085000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 193.195000 6.085000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 193.595000 6.085000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 193.995000 6.085000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 194.395000 6.085000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885000 194.795000 6.085000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 197.250000 50.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 197.650000 50.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 198.050000 50.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 198.450000 50.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 198.850000 50.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 199.250000 50.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.260000 199.650000 50.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 25.850000 50.740000 26.170000 ;
      LAYER met4 ;
        RECT 50.420000 25.850000 50.740000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 26.280000 50.740000 26.600000 ;
      LAYER met4 ;
        RECT 50.420000 26.280000 50.740000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 26.710000 50.740000 27.030000 ;
      LAYER met4 ;
        RECT 50.420000 26.710000 50.740000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 27.140000 50.740000 27.460000 ;
      LAYER met4 ;
        RECT 50.420000 27.140000 50.740000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 27.570000 50.740000 27.890000 ;
      LAYER met4 ;
        RECT 50.420000 27.570000 50.740000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 28.000000 50.740000 28.320000 ;
      LAYER met4 ;
        RECT 50.420000 28.000000 50.740000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 28.430000 50.740000 28.750000 ;
      LAYER met4 ;
        RECT 50.420000 28.430000 50.740000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 28.860000 50.740000 29.180000 ;
      LAYER met4 ;
        RECT 50.420000 28.860000 50.740000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 29.290000 50.740000 29.610000 ;
      LAYER met4 ;
        RECT 50.420000 29.290000 50.740000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 29.720000 50.740000 30.040000 ;
      LAYER met4 ;
        RECT 50.420000 29.720000 50.740000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 30.150000 50.740000 30.470000 ;
      LAYER met4 ;
        RECT 50.420000 30.150000 50.740000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 197.250000 50.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 197.650000 50.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 198.050000 50.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 198.450000 50.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 198.850000 50.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 199.250000 50.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 199.650000 50.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 25.850000 51.150000 26.170000 ;
      LAYER met4 ;
        RECT 50.830000 25.850000 51.150000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 26.280000 51.150000 26.600000 ;
      LAYER met4 ;
        RECT 50.830000 26.280000 51.150000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 26.710000 51.150000 27.030000 ;
      LAYER met4 ;
        RECT 50.830000 26.710000 51.150000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 27.140000 51.150000 27.460000 ;
      LAYER met4 ;
        RECT 50.830000 27.140000 51.150000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 27.570000 51.150000 27.890000 ;
      LAYER met4 ;
        RECT 50.830000 27.570000 51.150000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 28.000000 51.150000 28.320000 ;
      LAYER met4 ;
        RECT 50.830000 28.000000 51.150000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 28.430000 51.150000 28.750000 ;
      LAYER met4 ;
        RECT 50.830000 28.430000 51.150000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 28.860000 51.150000 29.180000 ;
      LAYER met4 ;
        RECT 50.830000 28.860000 51.150000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 29.290000 51.150000 29.610000 ;
      LAYER met4 ;
        RECT 50.830000 29.290000 51.150000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 29.720000 51.150000 30.040000 ;
      LAYER met4 ;
        RECT 50.830000 29.720000 51.150000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 30.150000 51.150000 30.470000 ;
      LAYER met4 ;
        RECT 50.830000 30.150000 51.150000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 197.250000 51.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 197.650000 51.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 198.050000 51.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 198.450000 51.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 198.850000 51.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 199.250000 51.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.060000 199.650000 51.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 25.850000 51.560000 26.170000 ;
      LAYER met4 ;
        RECT 51.240000 25.850000 51.560000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 26.280000 51.560000 26.600000 ;
      LAYER met4 ;
        RECT 51.240000 26.280000 51.560000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 26.710000 51.560000 27.030000 ;
      LAYER met4 ;
        RECT 51.240000 26.710000 51.560000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 27.140000 51.560000 27.460000 ;
      LAYER met4 ;
        RECT 51.240000 27.140000 51.560000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 27.570000 51.560000 27.890000 ;
      LAYER met4 ;
        RECT 51.240000 27.570000 51.560000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 28.000000 51.560000 28.320000 ;
      LAYER met4 ;
        RECT 51.240000 28.000000 51.560000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 28.430000 51.560000 28.750000 ;
      LAYER met4 ;
        RECT 51.240000 28.430000 51.560000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 28.860000 51.560000 29.180000 ;
      LAYER met4 ;
        RECT 51.240000 28.860000 51.560000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 29.290000 51.560000 29.610000 ;
      LAYER met4 ;
        RECT 51.240000 29.290000 51.560000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 29.720000 51.560000 30.040000 ;
      LAYER met4 ;
        RECT 51.240000 29.720000 51.560000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 30.150000 51.560000 30.470000 ;
      LAYER met4 ;
        RECT 51.240000 30.150000 51.560000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 197.250000 51.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 197.650000 51.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 198.050000 51.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 198.450000 51.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 198.850000 51.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 199.250000 51.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.460000 199.650000 51.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 25.850000 51.970000 26.170000 ;
      LAYER met4 ;
        RECT 51.650000 25.850000 51.970000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 26.280000 51.970000 26.600000 ;
      LAYER met4 ;
        RECT 51.650000 26.280000 51.970000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 26.710000 51.970000 27.030000 ;
      LAYER met4 ;
        RECT 51.650000 26.710000 51.970000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 27.140000 51.970000 27.460000 ;
      LAYER met4 ;
        RECT 51.650000 27.140000 51.970000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 27.570000 51.970000 27.890000 ;
      LAYER met4 ;
        RECT 51.650000 27.570000 51.970000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 28.000000 51.970000 28.320000 ;
      LAYER met4 ;
        RECT 51.650000 28.000000 51.970000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 28.430000 51.970000 28.750000 ;
      LAYER met4 ;
        RECT 51.650000 28.430000 51.970000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 28.860000 51.970000 29.180000 ;
      LAYER met4 ;
        RECT 51.650000 28.860000 51.970000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 29.290000 51.970000 29.610000 ;
      LAYER met4 ;
        RECT 51.650000 29.290000 51.970000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 29.720000 51.970000 30.040000 ;
      LAYER met4 ;
        RECT 51.650000 29.720000 51.970000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 30.150000 51.970000 30.470000 ;
      LAYER met4 ;
        RECT 51.650000 30.150000 51.970000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 197.250000 52.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 197.650000 52.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 198.050000 52.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 198.450000 52.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 198.850000 52.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 199.250000 52.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.860000 199.650000 52.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 25.850000 52.380000 26.170000 ;
      LAYER met4 ;
        RECT 52.060000 25.850000 52.380000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 26.280000 52.380000 26.600000 ;
      LAYER met4 ;
        RECT 52.060000 26.280000 52.380000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 26.710000 52.380000 27.030000 ;
      LAYER met4 ;
        RECT 52.060000 26.710000 52.380000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 27.140000 52.380000 27.460000 ;
      LAYER met4 ;
        RECT 52.060000 27.140000 52.380000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 27.570000 52.380000 27.890000 ;
      LAYER met4 ;
        RECT 52.060000 27.570000 52.380000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 28.000000 52.380000 28.320000 ;
      LAYER met4 ;
        RECT 52.060000 28.000000 52.380000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 28.430000 52.380000 28.750000 ;
      LAYER met4 ;
        RECT 52.060000 28.430000 52.380000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 28.860000 52.380000 29.180000 ;
      LAYER met4 ;
        RECT 52.060000 28.860000 52.380000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 29.290000 52.380000 29.610000 ;
      LAYER met4 ;
        RECT 52.060000 29.290000 52.380000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 29.720000 52.380000 30.040000 ;
      LAYER met4 ;
        RECT 52.060000 29.720000 52.380000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 30.150000 52.380000 30.470000 ;
      LAYER met4 ;
        RECT 52.060000 30.150000 52.380000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 197.250000 52.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 197.650000 52.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 198.050000 52.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 198.450000 52.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 198.850000 52.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 199.250000 52.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.260000 199.650000 52.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 25.850000 52.790000 26.170000 ;
      LAYER met4 ;
        RECT 52.470000 25.850000 52.790000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 26.280000 52.790000 26.600000 ;
      LAYER met4 ;
        RECT 52.470000 26.280000 52.790000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 26.710000 52.790000 27.030000 ;
      LAYER met4 ;
        RECT 52.470000 26.710000 52.790000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 27.140000 52.790000 27.460000 ;
      LAYER met4 ;
        RECT 52.470000 27.140000 52.790000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 27.570000 52.790000 27.890000 ;
      LAYER met4 ;
        RECT 52.470000 27.570000 52.790000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 28.000000 52.790000 28.320000 ;
      LAYER met4 ;
        RECT 52.470000 28.000000 52.790000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 28.430000 52.790000 28.750000 ;
      LAYER met4 ;
        RECT 52.470000 28.430000 52.790000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 28.860000 52.790000 29.180000 ;
      LAYER met4 ;
        RECT 52.470000 28.860000 52.790000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 29.290000 52.790000 29.610000 ;
      LAYER met4 ;
        RECT 52.470000 29.290000 52.790000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 29.720000 52.790000 30.040000 ;
      LAYER met4 ;
        RECT 52.470000 29.720000 52.790000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 30.150000 52.790000 30.470000 ;
      LAYER met4 ;
        RECT 52.470000 30.150000 52.790000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 197.250000 52.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 197.650000 52.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 198.050000 52.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 198.450000 52.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 198.850000 52.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 199.250000 52.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.660000 199.650000 52.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 25.850000 53.200000 26.170000 ;
      LAYER met4 ;
        RECT 52.880000 25.850000 53.200000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 26.280000 53.200000 26.600000 ;
      LAYER met4 ;
        RECT 52.880000 26.280000 53.200000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 26.710000 53.200000 27.030000 ;
      LAYER met4 ;
        RECT 52.880000 26.710000 53.200000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 27.140000 53.200000 27.460000 ;
      LAYER met4 ;
        RECT 52.880000 27.140000 53.200000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 27.570000 53.200000 27.890000 ;
      LAYER met4 ;
        RECT 52.880000 27.570000 53.200000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 28.000000 53.200000 28.320000 ;
      LAYER met4 ;
        RECT 52.880000 28.000000 53.200000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 28.430000 53.200000 28.750000 ;
      LAYER met4 ;
        RECT 52.880000 28.430000 53.200000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 28.860000 53.200000 29.180000 ;
      LAYER met4 ;
        RECT 52.880000 28.860000 53.200000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 29.290000 53.200000 29.610000 ;
      LAYER met4 ;
        RECT 52.880000 29.290000 53.200000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 29.720000 53.200000 30.040000 ;
      LAYER met4 ;
        RECT 52.880000 29.720000 53.200000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 30.150000 53.200000 30.470000 ;
      LAYER met4 ;
        RECT 52.880000 30.150000 53.200000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 197.250000 53.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 197.650000 53.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 198.050000 53.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 198.450000 53.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 198.850000 53.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 199.250000 53.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.060000 199.650000 53.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 25.850000 53.605000 26.170000 ;
      LAYER met4 ;
        RECT 53.285000 25.850000 53.605000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 26.280000 53.605000 26.600000 ;
      LAYER met4 ;
        RECT 53.285000 26.280000 53.605000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 26.710000 53.605000 27.030000 ;
      LAYER met4 ;
        RECT 53.285000 26.710000 53.605000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 27.140000 53.605000 27.460000 ;
      LAYER met4 ;
        RECT 53.285000 27.140000 53.605000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 27.570000 53.605000 27.890000 ;
      LAYER met4 ;
        RECT 53.285000 27.570000 53.605000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 28.000000 53.605000 28.320000 ;
      LAYER met4 ;
        RECT 53.285000 28.000000 53.605000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 28.430000 53.605000 28.750000 ;
      LAYER met4 ;
        RECT 53.285000 28.430000 53.605000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 28.860000 53.605000 29.180000 ;
      LAYER met4 ;
        RECT 53.285000 28.860000 53.605000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 29.290000 53.605000 29.610000 ;
      LAYER met4 ;
        RECT 53.285000 29.290000 53.605000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 29.720000 53.605000 30.040000 ;
      LAYER met4 ;
        RECT 53.285000 29.720000 53.605000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 30.150000 53.605000 30.470000 ;
      LAYER met4 ;
        RECT 53.285000 30.150000 53.605000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 197.250000 53.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 197.650000 53.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 198.050000 53.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 198.450000 53.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 198.850000 53.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 199.250000 53.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.460000 199.650000 53.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 25.850000 54.010000 26.170000 ;
      LAYER met4 ;
        RECT 53.690000 25.850000 54.010000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 26.280000 54.010000 26.600000 ;
      LAYER met4 ;
        RECT 53.690000 26.280000 54.010000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 26.710000 54.010000 27.030000 ;
      LAYER met4 ;
        RECT 53.690000 26.710000 54.010000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 27.140000 54.010000 27.460000 ;
      LAYER met4 ;
        RECT 53.690000 27.140000 54.010000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 27.570000 54.010000 27.890000 ;
      LAYER met4 ;
        RECT 53.690000 27.570000 54.010000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 28.000000 54.010000 28.320000 ;
      LAYER met4 ;
        RECT 53.690000 28.000000 54.010000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 28.430000 54.010000 28.750000 ;
      LAYER met4 ;
        RECT 53.690000 28.430000 54.010000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 28.860000 54.010000 29.180000 ;
      LAYER met4 ;
        RECT 53.690000 28.860000 54.010000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 29.290000 54.010000 29.610000 ;
      LAYER met4 ;
        RECT 53.690000 29.290000 54.010000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 29.720000 54.010000 30.040000 ;
      LAYER met4 ;
        RECT 53.690000 29.720000 54.010000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 30.150000 54.010000 30.470000 ;
      LAYER met4 ;
        RECT 53.690000 30.150000 54.010000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 197.250000 54.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 197.650000 54.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 198.050000 54.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 198.450000 54.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 198.850000 54.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 199.250000 54.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.860000 199.650000 54.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 25.850000 54.415000 26.170000 ;
      LAYER met4 ;
        RECT 54.095000 25.850000 54.415000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 26.280000 54.415000 26.600000 ;
      LAYER met4 ;
        RECT 54.095000 26.280000 54.415000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 26.710000 54.415000 27.030000 ;
      LAYER met4 ;
        RECT 54.095000 26.710000 54.415000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 27.140000 54.415000 27.460000 ;
      LAYER met4 ;
        RECT 54.095000 27.140000 54.415000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 27.570000 54.415000 27.890000 ;
      LAYER met4 ;
        RECT 54.095000 27.570000 54.415000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 28.000000 54.415000 28.320000 ;
      LAYER met4 ;
        RECT 54.095000 28.000000 54.415000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 28.430000 54.415000 28.750000 ;
      LAYER met4 ;
        RECT 54.095000 28.430000 54.415000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 28.860000 54.415000 29.180000 ;
      LAYER met4 ;
        RECT 54.095000 28.860000 54.415000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 29.290000 54.415000 29.610000 ;
      LAYER met4 ;
        RECT 54.095000 29.290000 54.415000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 29.720000 54.415000 30.040000 ;
      LAYER met4 ;
        RECT 54.095000 29.720000 54.415000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 30.150000 54.415000 30.470000 ;
      LAYER met4 ;
        RECT 54.095000 30.150000 54.415000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 197.250000 54.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 197.650000 54.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 198.050000 54.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 198.450000 54.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 198.850000 54.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 199.250000 54.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.260000 199.650000 54.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 25.850000 54.820000 26.170000 ;
      LAYER met4 ;
        RECT 54.500000 25.850000 54.820000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 26.280000 54.820000 26.600000 ;
      LAYER met4 ;
        RECT 54.500000 26.280000 54.820000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 26.710000 54.820000 27.030000 ;
      LAYER met4 ;
        RECT 54.500000 26.710000 54.820000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 27.140000 54.820000 27.460000 ;
      LAYER met4 ;
        RECT 54.500000 27.140000 54.820000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 27.570000 54.820000 27.890000 ;
      LAYER met4 ;
        RECT 54.500000 27.570000 54.820000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 28.000000 54.820000 28.320000 ;
      LAYER met4 ;
        RECT 54.500000 28.000000 54.820000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 28.430000 54.820000 28.750000 ;
      LAYER met4 ;
        RECT 54.500000 28.430000 54.820000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 28.860000 54.820000 29.180000 ;
      LAYER met4 ;
        RECT 54.500000 28.860000 54.820000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 29.290000 54.820000 29.610000 ;
      LAYER met4 ;
        RECT 54.500000 29.290000 54.820000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 29.720000 54.820000 30.040000 ;
      LAYER met4 ;
        RECT 54.500000 29.720000 54.820000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 30.150000 54.820000 30.470000 ;
      LAYER met4 ;
        RECT 54.500000 30.150000 54.820000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 197.250000 54.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 197.650000 54.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 198.050000 54.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 198.450000 54.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 198.850000 54.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 199.250000 54.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.660000 199.650000 54.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 25.850000 55.225000 26.170000 ;
      LAYER met4 ;
        RECT 54.905000 25.850000 55.225000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 26.280000 55.225000 26.600000 ;
      LAYER met4 ;
        RECT 54.905000 26.280000 55.225000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 26.710000 55.225000 27.030000 ;
      LAYER met4 ;
        RECT 54.905000 26.710000 55.225000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 27.140000 55.225000 27.460000 ;
      LAYER met4 ;
        RECT 54.905000 27.140000 55.225000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 27.570000 55.225000 27.890000 ;
      LAYER met4 ;
        RECT 54.905000 27.570000 55.225000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 28.000000 55.225000 28.320000 ;
      LAYER met4 ;
        RECT 54.905000 28.000000 55.225000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 28.430000 55.225000 28.750000 ;
      LAYER met4 ;
        RECT 54.905000 28.430000 55.225000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 28.860000 55.225000 29.180000 ;
      LAYER met4 ;
        RECT 54.905000 28.860000 55.225000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 29.290000 55.225000 29.610000 ;
      LAYER met4 ;
        RECT 54.905000 29.290000 55.225000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 29.720000 55.225000 30.040000 ;
      LAYER met4 ;
        RECT 54.905000 29.720000 55.225000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 30.150000 55.225000 30.470000 ;
      LAYER met4 ;
        RECT 54.905000 30.150000 55.225000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 197.250000 55.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 197.650000 55.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 198.050000 55.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 198.450000 55.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 198.850000 55.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 199.250000 55.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.060000 199.650000 55.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 25.850000 55.630000 26.170000 ;
      LAYER met4 ;
        RECT 55.310000 25.850000 55.630000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 26.280000 55.630000 26.600000 ;
      LAYER met4 ;
        RECT 55.310000 26.280000 55.630000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 26.710000 55.630000 27.030000 ;
      LAYER met4 ;
        RECT 55.310000 26.710000 55.630000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 27.140000 55.630000 27.460000 ;
      LAYER met4 ;
        RECT 55.310000 27.140000 55.630000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 27.570000 55.630000 27.890000 ;
      LAYER met4 ;
        RECT 55.310000 27.570000 55.630000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 28.000000 55.630000 28.320000 ;
      LAYER met4 ;
        RECT 55.310000 28.000000 55.630000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 28.430000 55.630000 28.750000 ;
      LAYER met4 ;
        RECT 55.310000 28.430000 55.630000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 28.860000 55.630000 29.180000 ;
      LAYER met4 ;
        RECT 55.310000 28.860000 55.630000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 29.290000 55.630000 29.610000 ;
      LAYER met4 ;
        RECT 55.310000 29.290000 55.630000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 29.720000 55.630000 30.040000 ;
      LAYER met4 ;
        RECT 55.310000 29.720000 55.630000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 30.150000 55.630000 30.470000 ;
      LAYER met4 ;
        RECT 55.310000 30.150000 55.630000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 197.250000 55.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 197.650000 55.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 198.050000 55.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 198.450000 55.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 198.850000 55.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 199.250000 55.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.460000 199.650000 55.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 25.850000 56.035000 26.170000 ;
      LAYER met4 ;
        RECT 55.715000 25.850000 56.035000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 26.280000 56.035000 26.600000 ;
      LAYER met4 ;
        RECT 55.715000 26.280000 56.035000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 26.710000 56.035000 27.030000 ;
      LAYER met4 ;
        RECT 55.715000 26.710000 56.035000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 27.140000 56.035000 27.460000 ;
      LAYER met4 ;
        RECT 55.715000 27.140000 56.035000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 27.570000 56.035000 27.890000 ;
      LAYER met4 ;
        RECT 55.715000 27.570000 56.035000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 28.000000 56.035000 28.320000 ;
      LAYER met4 ;
        RECT 55.715000 28.000000 56.035000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 28.430000 56.035000 28.750000 ;
      LAYER met4 ;
        RECT 55.715000 28.430000 56.035000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 28.860000 56.035000 29.180000 ;
      LAYER met4 ;
        RECT 55.715000 28.860000 56.035000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 29.290000 56.035000 29.610000 ;
      LAYER met4 ;
        RECT 55.715000 29.290000 56.035000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 29.720000 56.035000 30.040000 ;
      LAYER met4 ;
        RECT 55.715000 29.720000 56.035000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 30.150000 56.035000 30.470000 ;
      LAYER met4 ;
        RECT 55.715000 30.150000 56.035000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 197.250000 56.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 197.650000 56.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 198.050000 56.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 198.450000 56.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 198.850000 56.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 199.250000 56.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.860000 199.650000 56.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 25.850000 56.440000 26.170000 ;
      LAYER met4 ;
        RECT 56.120000 25.850000 56.440000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 26.280000 56.440000 26.600000 ;
      LAYER met4 ;
        RECT 56.120000 26.280000 56.440000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 26.710000 56.440000 27.030000 ;
      LAYER met4 ;
        RECT 56.120000 26.710000 56.440000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 27.140000 56.440000 27.460000 ;
      LAYER met4 ;
        RECT 56.120000 27.140000 56.440000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 27.570000 56.440000 27.890000 ;
      LAYER met4 ;
        RECT 56.120000 27.570000 56.440000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 28.000000 56.440000 28.320000 ;
      LAYER met4 ;
        RECT 56.120000 28.000000 56.440000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 28.430000 56.440000 28.750000 ;
      LAYER met4 ;
        RECT 56.120000 28.430000 56.440000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 28.860000 56.440000 29.180000 ;
      LAYER met4 ;
        RECT 56.120000 28.860000 56.440000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 29.290000 56.440000 29.610000 ;
      LAYER met4 ;
        RECT 56.120000 29.290000 56.440000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 29.720000 56.440000 30.040000 ;
      LAYER met4 ;
        RECT 56.120000 29.720000 56.440000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 30.150000 56.440000 30.470000 ;
      LAYER met4 ;
        RECT 56.120000 30.150000 56.440000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 197.250000 56.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 197.650000 56.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 198.050000 56.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 198.450000 56.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 198.850000 56.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 199.250000 56.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260000 199.650000 56.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 25.850000 56.845000 26.170000 ;
      LAYER met4 ;
        RECT 56.525000 25.850000 56.845000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 26.280000 56.845000 26.600000 ;
      LAYER met4 ;
        RECT 56.525000 26.280000 56.845000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 26.710000 56.845000 27.030000 ;
      LAYER met4 ;
        RECT 56.525000 26.710000 56.845000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 27.140000 56.845000 27.460000 ;
      LAYER met4 ;
        RECT 56.525000 27.140000 56.845000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 27.570000 56.845000 27.890000 ;
      LAYER met4 ;
        RECT 56.525000 27.570000 56.845000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 28.000000 56.845000 28.320000 ;
      LAYER met4 ;
        RECT 56.525000 28.000000 56.845000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 28.430000 56.845000 28.750000 ;
      LAYER met4 ;
        RECT 56.525000 28.430000 56.845000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 28.860000 56.845000 29.180000 ;
      LAYER met4 ;
        RECT 56.525000 28.860000 56.845000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 29.290000 56.845000 29.610000 ;
      LAYER met4 ;
        RECT 56.525000 29.290000 56.845000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 29.720000 56.845000 30.040000 ;
      LAYER met4 ;
        RECT 56.525000 29.720000 56.845000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 30.150000 56.845000 30.470000 ;
      LAYER met4 ;
        RECT 56.525000 30.150000 56.845000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 197.250000 56.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 197.650000 56.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 198.050000 56.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 198.450000 56.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 198.850000 56.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 199.250000 56.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.660000 199.650000 56.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 25.850000 57.250000 26.170000 ;
      LAYER met4 ;
        RECT 56.930000 25.850000 57.250000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 26.280000 57.250000 26.600000 ;
      LAYER met4 ;
        RECT 56.930000 26.280000 57.250000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 26.710000 57.250000 27.030000 ;
      LAYER met4 ;
        RECT 56.930000 26.710000 57.250000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 27.140000 57.250000 27.460000 ;
      LAYER met4 ;
        RECT 56.930000 27.140000 57.250000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 27.570000 57.250000 27.890000 ;
      LAYER met4 ;
        RECT 56.930000 27.570000 57.250000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 28.000000 57.250000 28.320000 ;
      LAYER met4 ;
        RECT 56.930000 28.000000 57.250000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 28.430000 57.250000 28.750000 ;
      LAYER met4 ;
        RECT 56.930000 28.430000 57.250000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 28.860000 57.250000 29.180000 ;
      LAYER met4 ;
        RECT 56.930000 28.860000 57.250000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 29.290000 57.250000 29.610000 ;
      LAYER met4 ;
        RECT 56.930000 29.290000 57.250000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 29.720000 57.250000 30.040000 ;
      LAYER met4 ;
        RECT 56.930000 29.720000 57.250000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 30.150000 57.250000 30.470000 ;
      LAYER met4 ;
        RECT 56.930000 30.150000 57.250000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 197.250000 57.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 197.650000 57.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 198.050000 57.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 198.450000 57.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 198.850000 57.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 199.250000 57.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.060000 199.650000 57.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 25.850000 57.655000 26.170000 ;
      LAYER met4 ;
        RECT 57.335000 25.850000 57.655000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 26.280000 57.655000 26.600000 ;
      LAYER met4 ;
        RECT 57.335000 26.280000 57.655000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 26.710000 57.655000 27.030000 ;
      LAYER met4 ;
        RECT 57.335000 26.710000 57.655000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 27.140000 57.655000 27.460000 ;
      LAYER met4 ;
        RECT 57.335000 27.140000 57.655000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 27.570000 57.655000 27.890000 ;
      LAYER met4 ;
        RECT 57.335000 27.570000 57.655000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 28.000000 57.655000 28.320000 ;
      LAYER met4 ;
        RECT 57.335000 28.000000 57.655000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 28.430000 57.655000 28.750000 ;
      LAYER met4 ;
        RECT 57.335000 28.430000 57.655000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 28.860000 57.655000 29.180000 ;
      LAYER met4 ;
        RECT 57.335000 28.860000 57.655000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 29.290000 57.655000 29.610000 ;
      LAYER met4 ;
        RECT 57.335000 29.290000 57.655000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 29.720000 57.655000 30.040000 ;
      LAYER met4 ;
        RECT 57.335000 29.720000 57.655000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 30.150000 57.655000 30.470000 ;
      LAYER met4 ;
        RECT 57.335000 30.150000 57.655000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 197.250000 57.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 197.650000 57.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 198.050000 57.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 198.450000 57.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 198.850000 57.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 199.250000 57.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.460000 199.650000 57.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 25.850000 58.060000 26.170000 ;
      LAYER met4 ;
        RECT 57.740000 25.850000 58.060000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 26.280000 58.060000 26.600000 ;
      LAYER met4 ;
        RECT 57.740000 26.280000 58.060000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 26.710000 58.060000 27.030000 ;
      LAYER met4 ;
        RECT 57.740000 26.710000 58.060000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 27.140000 58.060000 27.460000 ;
      LAYER met4 ;
        RECT 57.740000 27.140000 58.060000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 27.570000 58.060000 27.890000 ;
      LAYER met4 ;
        RECT 57.740000 27.570000 58.060000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 28.000000 58.060000 28.320000 ;
      LAYER met4 ;
        RECT 57.740000 28.000000 58.060000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 28.430000 58.060000 28.750000 ;
      LAYER met4 ;
        RECT 57.740000 28.430000 58.060000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 28.860000 58.060000 29.180000 ;
      LAYER met4 ;
        RECT 57.740000 28.860000 58.060000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 29.290000 58.060000 29.610000 ;
      LAYER met4 ;
        RECT 57.740000 29.290000 58.060000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 29.720000 58.060000 30.040000 ;
      LAYER met4 ;
        RECT 57.740000 29.720000 58.060000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 30.150000 58.060000 30.470000 ;
      LAYER met4 ;
        RECT 57.740000 30.150000 58.060000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 197.250000 58.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 197.650000 58.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 198.050000 58.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 198.450000 58.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 198.850000 58.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 199.250000 58.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.860000 199.650000 58.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 25.850000 58.465000 26.170000 ;
      LAYER met4 ;
        RECT 58.145000 25.850000 58.465000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 26.280000 58.465000 26.600000 ;
      LAYER met4 ;
        RECT 58.145000 26.280000 58.465000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 26.710000 58.465000 27.030000 ;
      LAYER met4 ;
        RECT 58.145000 26.710000 58.465000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 27.140000 58.465000 27.460000 ;
      LAYER met4 ;
        RECT 58.145000 27.140000 58.465000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 27.570000 58.465000 27.890000 ;
      LAYER met4 ;
        RECT 58.145000 27.570000 58.465000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 28.000000 58.465000 28.320000 ;
      LAYER met4 ;
        RECT 58.145000 28.000000 58.465000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 28.430000 58.465000 28.750000 ;
      LAYER met4 ;
        RECT 58.145000 28.430000 58.465000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 28.860000 58.465000 29.180000 ;
      LAYER met4 ;
        RECT 58.145000 28.860000 58.465000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 29.290000 58.465000 29.610000 ;
      LAYER met4 ;
        RECT 58.145000 29.290000 58.465000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 29.720000 58.465000 30.040000 ;
      LAYER met4 ;
        RECT 58.145000 29.720000 58.465000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 30.150000 58.465000 30.470000 ;
      LAYER met4 ;
        RECT 58.145000 30.150000 58.465000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 197.250000 58.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 197.650000 58.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 198.050000 58.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 198.450000 58.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 198.850000 58.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 199.250000 58.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.260000 199.650000 58.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 25.850000 58.870000 26.170000 ;
      LAYER met4 ;
        RECT 58.550000 25.850000 58.870000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 26.280000 58.870000 26.600000 ;
      LAYER met4 ;
        RECT 58.550000 26.280000 58.870000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 26.710000 58.870000 27.030000 ;
      LAYER met4 ;
        RECT 58.550000 26.710000 58.870000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 27.140000 58.870000 27.460000 ;
      LAYER met4 ;
        RECT 58.550000 27.140000 58.870000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 27.570000 58.870000 27.890000 ;
      LAYER met4 ;
        RECT 58.550000 27.570000 58.870000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 28.000000 58.870000 28.320000 ;
      LAYER met4 ;
        RECT 58.550000 28.000000 58.870000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 28.430000 58.870000 28.750000 ;
      LAYER met4 ;
        RECT 58.550000 28.430000 58.870000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 28.860000 58.870000 29.180000 ;
      LAYER met4 ;
        RECT 58.550000 28.860000 58.870000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 29.290000 58.870000 29.610000 ;
      LAYER met4 ;
        RECT 58.550000 29.290000 58.870000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 29.720000 58.870000 30.040000 ;
      LAYER met4 ;
        RECT 58.550000 29.720000 58.870000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 30.150000 58.870000 30.470000 ;
      LAYER met4 ;
        RECT 58.550000 30.150000 58.870000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 197.250000 58.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 197.650000 58.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 198.050000 58.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 198.450000 58.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 198.850000 58.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 199.250000 58.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.660000 199.650000 58.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 25.850000 59.275000 26.170000 ;
      LAYER met4 ;
        RECT 58.955000 25.850000 59.275000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 26.280000 59.275000 26.600000 ;
      LAYER met4 ;
        RECT 58.955000 26.280000 59.275000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 26.710000 59.275000 27.030000 ;
      LAYER met4 ;
        RECT 58.955000 26.710000 59.275000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 27.140000 59.275000 27.460000 ;
      LAYER met4 ;
        RECT 58.955000 27.140000 59.275000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 27.570000 59.275000 27.890000 ;
      LAYER met4 ;
        RECT 58.955000 27.570000 59.275000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 28.000000 59.275000 28.320000 ;
      LAYER met4 ;
        RECT 58.955000 28.000000 59.275000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 28.430000 59.275000 28.750000 ;
      LAYER met4 ;
        RECT 58.955000 28.430000 59.275000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 28.860000 59.275000 29.180000 ;
      LAYER met4 ;
        RECT 58.955000 28.860000 59.275000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 29.290000 59.275000 29.610000 ;
      LAYER met4 ;
        RECT 58.955000 29.290000 59.275000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 29.720000 59.275000 30.040000 ;
      LAYER met4 ;
        RECT 58.955000 29.720000 59.275000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 30.150000 59.275000 30.470000 ;
      LAYER met4 ;
        RECT 58.955000 30.150000 59.275000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 197.250000 59.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 197.650000 59.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 198.050000 59.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 198.450000 59.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 198.850000 59.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 199.250000 59.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.060000 199.650000 59.260000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 25.850000 59.680000 26.170000 ;
      LAYER met4 ;
        RECT 59.360000 25.850000 59.680000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 26.280000 59.680000 26.600000 ;
      LAYER met4 ;
        RECT 59.360000 26.280000 59.680000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 26.710000 59.680000 27.030000 ;
      LAYER met4 ;
        RECT 59.360000 26.710000 59.680000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 27.140000 59.680000 27.460000 ;
      LAYER met4 ;
        RECT 59.360000 27.140000 59.680000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 27.570000 59.680000 27.890000 ;
      LAYER met4 ;
        RECT 59.360000 27.570000 59.680000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 28.000000 59.680000 28.320000 ;
      LAYER met4 ;
        RECT 59.360000 28.000000 59.680000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 28.430000 59.680000 28.750000 ;
      LAYER met4 ;
        RECT 59.360000 28.430000 59.680000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 28.860000 59.680000 29.180000 ;
      LAYER met4 ;
        RECT 59.360000 28.860000 59.680000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 29.290000 59.680000 29.610000 ;
      LAYER met4 ;
        RECT 59.360000 29.290000 59.680000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 29.720000 59.680000 30.040000 ;
      LAYER met4 ;
        RECT 59.360000 29.720000 59.680000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 30.150000 59.680000 30.470000 ;
      LAYER met4 ;
        RECT 59.360000 30.150000 59.680000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 197.250000 59.660000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 197.650000 59.660000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 198.050000 59.660000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 198.450000 59.660000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 198.850000 59.660000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 199.250000 59.660000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.460000 199.650000 59.660000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 25.850000 60.085000 26.170000 ;
      LAYER met4 ;
        RECT 59.765000 25.850000 60.085000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 26.280000 60.085000 26.600000 ;
      LAYER met4 ;
        RECT 59.765000 26.280000 60.085000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 26.710000 60.085000 27.030000 ;
      LAYER met4 ;
        RECT 59.765000 26.710000 60.085000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 27.140000 60.085000 27.460000 ;
      LAYER met4 ;
        RECT 59.765000 27.140000 60.085000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 27.570000 60.085000 27.890000 ;
      LAYER met4 ;
        RECT 59.765000 27.570000 60.085000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 28.000000 60.085000 28.320000 ;
      LAYER met4 ;
        RECT 59.765000 28.000000 60.085000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 28.430000 60.085000 28.750000 ;
      LAYER met4 ;
        RECT 59.765000 28.430000 60.085000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 28.860000 60.085000 29.180000 ;
      LAYER met4 ;
        RECT 59.765000 28.860000 60.085000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 29.290000 60.085000 29.610000 ;
      LAYER met4 ;
        RECT 59.765000 29.290000 60.085000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 29.720000 60.085000 30.040000 ;
      LAYER met4 ;
        RECT 59.765000 29.720000 60.085000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 30.150000 60.085000 30.470000 ;
      LAYER met4 ;
        RECT 59.765000 30.150000 60.085000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 197.250000 60.060000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 197.650000 60.060000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 198.050000 60.060000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 198.450000 60.060000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 198.850000 60.060000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 199.250000 60.060000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.860000 199.650000 60.060000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 195.140000 6.545000 195.460000 ;
      LAYER met4 ;
        RECT 6.225000 195.140000 6.545000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 195.545000 6.545000 195.865000 ;
      LAYER met4 ;
        RECT 6.225000 195.545000 6.545000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 195.950000 6.545000 196.270000 ;
      LAYER met4 ;
        RECT 6.225000 195.950000 6.545000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 196.355000 6.545000 196.675000 ;
      LAYER met4 ;
        RECT 6.225000 196.355000 6.545000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 196.760000 6.545000 197.080000 ;
      LAYER met4 ;
        RECT 6.225000 196.760000 6.545000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 197.165000 6.545000 197.485000 ;
      LAYER met4 ;
        RECT 6.225000 197.165000 6.545000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 197.570000 6.545000 197.890000 ;
      LAYER met4 ;
        RECT 6.225000 197.570000 6.545000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 197.975000 6.545000 198.295000 ;
      LAYER met4 ;
        RECT 6.225000 197.975000 6.545000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 198.380000 6.545000 198.700000 ;
      LAYER met4 ;
        RECT 6.225000 198.380000 6.545000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 198.785000 6.545000 199.105000 ;
      LAYER met4 ;
        RECT 6.225000 198.785000 6.545000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 199.190000 6.545000 199.510000 ;
      LAYER met4 ;
        RECT 6.225000 199.190000 6.545000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 199.595000 6.545000 199.915000 ;
      LAYER met4 ;
        RECT 6.225000 199.595000 6.545000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 25.850000 6.545000 26.170000 ;
      LAYER met4 ;
        RECT 6.225000 25.850000 6.545000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 26.280000 6.545000 26.600000 ;
      LAYER met4 ;
        RECT 6.225000 26.280000 6.545000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 26.710000 6.545000 27.030000 ;
      LAYER met4 ;
        RECT 6.225000 26.710000 6.545000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 27.140000 6.545000 27.460000 ;
      LAYER met4 ;
        RECT 6.225000 27.140000 6.545000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 27.570000 6.545000 27.890000 ;
      LAYER met4 ;
        RECT 6.225000 27.570000 6.545000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 28.000000 6.545000 28.320000 ;
      LAYER met4 ;
        RECT 6.225000 28.000000 6.545000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 28.430000 6.545000 28.750000 ;
      LAYER met4 ;
        RECT 6.225000 28.430000 6.545000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 28.860000 6.545000 29.180000 ;
      LAYER met4 ;
        RECT 6.225000 28.860000 6.545000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 29.290000 6.545000 29.610000 ;
      LAYER met4 ;
        RECT 6.225000 29.290000 6.545000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 29.720000 6.545000 30.040000 ;
      LAYER met4 ;
        RECT 6.225000 29.720000 6.545000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 30.150000 6.545000 30.470000 ;
      LAYER met4 ;
        RECT 6.225000 30.150000 6.545000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 175.995000 6.485000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 176.395000 6.485000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 176.795000 6.485000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 177.195000 6.485000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 177.595000 6.485000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 177.995000 6.485000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 178.395000 6.485000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 178.795000 6.485000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 179.195000 6.485000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 179.595000 6.485000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 179.995000 6.485000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 180.395000 6.485000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 180.795000 6.485000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 181.195000 6.485000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 181.595000 6.485000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 181.995000 6.485000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 182.395000 6.485000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 182.795000 6.485000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 183.195000 6.485000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 183.595000 6.485000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 183.995000 6.485000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 184.395000 6.485000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 184.795000 6.485000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 185.195000 6.485000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 185.595000 6.485000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 185.995000 6.485000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 186.395000 6.485000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 186.795000 6.485000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 187.195000 6.485000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 187.595000 6.485000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 187.995000 6.485000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 188.395000 6.485000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 188.795000 6.485000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 189.195000 6.485000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 189.595000 6.485000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 189.995000 6.485000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 190.395000 6.485000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 190.795000 6.485000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 191.195000 6.485000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 191.595000 6.485000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 191.995000 6.485000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 192.395000 6.485000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 192.795000 6.485000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 193.195000 6.485000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 193.595000 6.485000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 193.995000 6.485000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 194.395000 6.485000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285000 194.795000 6.485000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 195.140000 6.945000 195.460000 ;
      LAYER met4 ;
        RECT 6.625000 195.140000 6.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 195.545000 6.945000 195.865000 ;
      LAYER met4 ;
        RECT 6.625000 195.545000 6.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 195.950000 6.945000 196.270000 ;
      LAYER met4 ;
        RECT 6.625000 195.950000 6.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 196.355000 6.945000 196.675000 ;
      LAYER met4 ;
        RECT 6.625000 196.355000 6.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 196.760000 6.945000 197.080000 ;
      LAYER met4 ;
        RECT 6.625000 196.760000 6.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 197.165000 6.945000 197.485000 ;
      LAYER met4 ;
        RECT 6.625000 197.165000 6.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 197.570000 6.945000 197.890000 ;
      LAYER met4 ;
        RECT 6.625000 197.570000 6.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 197.975000 6.945000 198.295000 ;
      LAYER met4 ;
        RECT 6.625000 197.975000 6.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 198.380000 6.945000 198.700000 ;
      LAYER met4 ;
        RECT 6.625000 198.380000 6.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 198.785000 6.945000 199.105000 ;
      LAYER met4 ;
        RECT 6.625000 198.785000 6.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 199.190000 6.945000 199.510000 ;
      LAYER met4 ;
        RECT 6.625000 199.190000 6.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625000 199.595000 6.945000 199.915000 ;
      LAYER met4 ;
        RECT 6.625000 199.595000 6.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 25.850000 6.950000 26.170000 ;
      LAYER met4 ;
        RECT 6.630000 25.850000 6.950000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 26.280000 6.950000 26.600000 ;
      LAYER met4 ;
        RECT 6.630000 26.280000 6.950000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 26.710000 6.950000 27.030000 ;
      LAYER met4 ;
        RECT 6.630000 26.710000 6.950000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 27.140000 6.950000 27.460000 ;
      LAYER met4 ;
        RECT 6.630000 27.140000 6.950000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 27.570000 6.950000 27.890000 ;
      LAYER met4 ;
        RECT 6.630000 27.570000 6.950000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 28.000000 6.950000 28.320000 ;
      LAYER met4 ;
        RECT 6.630000 28.000000 6.950000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 28.430000 6.950000 28.750000 ;
      LAYER met4 ;
        RECT 6.630000 28.430000 6.950000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 28.860000 6.950000 29.180000 ;
      LAYER met4 ;
        RECT 6.630000 28.860000 6.950000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 29.290000 6.950000 29.610000 ;
      LAYER met4 ;
        RECT 6.630000 29.290000 6.950000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 29.720000 6.950000 30.040000 ;
      LAYER met4 ;
        RECT 6.630000 29.720000 6.950000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 30.150000 6.950000 30.470000 ;
      LAYER met4 ;
        RECT 6.630000 30.150000 6.950000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 175.995000 6.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 176.395000 6.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 176.795000 6.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 177.195000 6.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 177.595000 6.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 177.995000 6.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 178.395000 6.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 178.795000 6.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 179.195000 6.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 179.595000 6.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 179.995000 6.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 180.395000 6.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 180.795000 6.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 181.195000 6.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 181.595000 6.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 181.995000 6.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 182.395000 6.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 182.795000 6.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 183.195000 6.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 183.595000 6.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 183.995000 6.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 184.395000 6.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 184.795000 6.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 185.195000 6.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 185.595000 6.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 185.995000 6.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 186.395000 6.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 186.795000 6.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 187.195000 6.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 187.595000 6.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 187.995000 6.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 188.395000 6.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 188.795000 6.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 189.195000 6.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 189.595000 6.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 189.995000 6.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 190.395000 6.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 190.795000 6.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 191.195000 6.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 191.595000 6.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 191.995000 6.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 192.395000 6.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 192.795000 6.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 193.195000 6.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 193.595000 6.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 193.995000 6.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 194.395000 6.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.685000 194.795000 6.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 25.850000 60.490000 26.170000 ;
      LAYER met4 ;
        RECT 60.170000 25.850000 60.490000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 26.280000 60.490000 26.600000 ;
      LAYER met4 ;
        RECT 60.170000 26.280000 60.490000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 26.710000 60.490000 27.030000 ;
      LAYER met4 ;
        RECT 60.170000 26.710000 60.490000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 27.140000 60.490000 27.460000 ;
      LAYER met4 ;
        RECT 60.170000 27.140000 60.490000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 27.570000 60.490000 27.890000 ;
      LAYER met4 ;
        RECT 60.170000 27.570000 60.490000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 28.000000 60.490000 28.320000 ;
      LAYER met4 ;
        RECT 60.170000 28.000000 60.490000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 28.430000 60.490000 28.750000 ;
      LAYER met4 ;
        RECT 60.170000 28.430000 60.490000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 28.860000 60.490000 29.180000 ;
      LAYER met4 ;
        RECT 60.170000 28.860000 60.490000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 29.290000 60.490000 29.610000 ;
      LAYER met4 ;
        RECT 60.170000 29.290000 60.490000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 29.720000 60.490000 30.040000 ;
      LAYER met4 ;
        RECT 60.170000 29.720000 60.490000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 30.150000 60.490000 30.470000 ;
      LAYER met4 ;
        RECT 60.170000 30.150000 60.490000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 197.250000 60.460000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 197.650000 60.460000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 198.050000 60.460000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 198.450000 60.460000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 198.850000 60.460000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 199.250000 60.460000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.260000 199.650000 60.460000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 25.850000 60.895000 26.170000 ;
      LAYER met4 ;
        RECT 60.575000 25.850000 60.895000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 26.280000 60.895000 26.600000 ;
      LAYER met4 ;
        RECT 60.575000 26.280000 60.895000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 26.710000 60.895000 27.030000 ;
      LAYER met4 ;
        RECT 60.575000 26.710000 60.895000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 27.140000 60.895000 27.460000 ;
      LAYER met4 ;
        RECT 60.575000 27.140000 60.895000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 27.570000 60.895000 27.890000 ;
      LAYER met4 ;
        RECT 60.575000 27.570000 60.895000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 28.000000 60.895000 28.320000 ;
      LAYER met4 ;
        RECT 60.575000 28.000000 60.895000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 28.430000 60.895000 28.750000 ;
      LAYER met4 ;
        RECT 60.575000 28.430000 60.895000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 28.860000 60.895000 29.180000 ;
      LAYER met4 ;
        RECT 60.575000 28.860000 60.895000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 29.290000 60.895000 29.610000 ;
      LAYER met4 ;
        RECT 60.575000 29.290000 60.895000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 29.720000 60.895000 30.040000 ;
      LAYER met4 ;
        RECT 60.575000 29.720000 60.895000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 30.150000 60.895000 30.470000 ;
      LAYER met4 ;
        RECT 60.575000 30.150000 60.895000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 197.250000 60.860000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 197.650000 60.860000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 198.050000 60.860000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 198.450000 60.860000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 198.850000 60.860000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 199.250000 60.860000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.660000 199.650000 60.860000 199.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.850000 196.235000 61.170000 196.555000 ;
      LAYER met4 ;
        RECT 60.850000 196.235000 61.170000 196.555000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.850000 196.645000 61.170000 196.965000 ;
      LAYER met4 ;
        RECT 60.850000 196.645000 61.170000 196.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 25.850000 61.300000 26.170000 ;
      LAYER met4 ;
        RECT 60.980000 25.850000 61.300000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 26.280000 61.300000 26.600000 ;
      LAYER met4 ;
        RECT 60.980000 26.280000 61.300000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 26.710000 61.300000 27.030000 ;
      LAYER met4 ;
        RECT 60.980000 26.710000 61.300000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 27.140000 61.300000 27.460000 ;
      LAYER met4 ;
        RECT 60.980000 27.140000 61.300000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 27.570000 61.300000 27.890000 ;
      LAYER met4 ;
        RECT 60.980000 27.570000 61.300000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 28.000000 61.300000 28.320000 ;
      LAYER met4 ;
        RECT 60.980000 28.000000 61.300000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 28.430000 61.300000 28.750000 ;
      LAYER met4 ;
        RECT 60.980000 28.430000 61.300000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 28.860000 61.300000 29.180000 ;
      LAYER met4 ;
        RECT 60.980000 28.860000 61.300000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 29.290000 61.300000 29.610000 ;
      LAYER met4 ;
        RECT 60.980000 29.290000 61.300000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 29.720000 61.300000 30.040000 ;
      LAYER met4 ;
        RECT 60.980000 29.720000 61.300000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 30.150000 61.300000 30.470000 ;
      LAYER met4 ;
        RECT 60.980000 30.150000 61.300000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.060000 197.250000 61.260000 197.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.060000 197.650000 61.260000 197.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.060000 198.050000 61.260000 198.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.060000 198.450000 61.260000 198.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.060000 198.850000 61.260000 199.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.060000 199.250000 61.260000 199.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 25.850000 61.705000 26.170000 ;
      LAYER met4 ;
        RECT 61.385000 25.850000 61.705000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 26.280000 61.705000 26.600000 ;
      LAYER met4 ;
        RECT 61.385000 26.280000 61.705000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 26.710000 61.705000 27.030000 ;
      LAYER met4 ;
        RECT 61.385000 26.710000 61.705000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 27.140000 61.705000 27.460000 ;
      LAYER met4 ;
        RECT 61.385000 27.140000 61.705000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 27.570000 61.705000 27.890000 ;
      LAYER met4 ;
        RECT 61.385000 27.570000 61.705000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 28.000000 61.705000 28.320000 ;
      LAYER met4 ;
        RECT 61.385000 28.000000 61.705000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 28.430000 61.705000 28.750000 ;
      LAYER met4 ;
        RECT 61.385000 28.430000 61.705000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 28.860000 61.705000 29.180000 ;
      LAYER met4 ;
        RECT 61.385000 28.860000 61.705000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 29.290000 61.705000 29.610000 ;
      LAYER met4 ;
        RECT 61.385000 29.290000 61.705000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 29.720000 61.705000 30.040000 ;
      LAYER met4 ;
        RECT 61.385000 29.720000 61.705000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 30.150000 61.705000 30.470000 ;
      LAYER met4 ;
        RECT 61.385000 30.150000 61.705000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 175.935000 74.250000 195.055000 ;
      LAYER met4 ;
        RECT 61.530000 175.935000 74.250000 195.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 195.140000 61.850000 195.460000 ;
      LAYER met4 ;
        RECT 61.530000 195.140000 61.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 195.545000 61.850000 195.865000 ;
      LAYER met4 ;
        RECT 61.530000 195.545000 61.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 195.950000 61.850000 196.270000 ;
      LAYER met4 ;
        RECT 61.530000 195.950000 61.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 196.355000 61.850000 196.675000 ;
      LAYER met4 ;
        RECT 61.530000 196.355000 61.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 196.760000 61.850000 197.080000 ;
      LAYER met4 ;
        RECT 61.530000 196.760000 61.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 197.165000 61.850000 197.485000 ;
      LAYER met4 ;
        RECT 61.530000 197.165000 61.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 197.570000 61.850000 197.890000 ;
      LAYER met4 ;
        RECT 61.530000 197.570000 61.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 197.975000 61.850000 198.295000 ;
      LAYER met4 ;
        RECT 61.530000 197.975000 61.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 198.380000 61.850000 198.700000 ;
      LAYER met4 ;
        RECT 61.530000 198.380000 61.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 198.785000 61.850000 199.105000 ;
      LAYER met4 ;
        RECT 61.530000 198.785000 61.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 199.190000 61.850000 199.510000 ;
      LAYER met4 ;
        RECT 61.530000 199.190000 61.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530000 199.595000 61.850000 199.915000 ;
      LAYER met4 ;
        RECT 61.530000 199.595000 61.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 175.995000 61.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 176.395000 61.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 176.795000 61.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 177.195000 61.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 177.595000 61.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 177.995000 61.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 178.395000 61.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 178.795000 61.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 179.195000 61.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 179.595000 61.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 179.995000 61.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 180.395000 61.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 180.795000 61.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 181.195000 61.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 181.595000 61.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 181.995000 61.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 182.395000 61.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 182.795000 61.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 183.195000 61.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 183.595000 61.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 183.995000 61.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 184.395000 61.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 184.795000 61.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 185.195000 61.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 185.595000 61.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 185.995000 61.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 186.395000 61.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 186.795000 61.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 187.195000 61.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 187.595000 61.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 187.995000 61.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 188.395000 61.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 188.795000 61.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 189.195000 61.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 189.595000 61.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 189.995000 61.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 190.395000 61.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 190.795000 61.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 191.195000 61.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 191.595000 61.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 191.995000 61.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 192.395000 61.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 192.795000 61.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 193.195000 61.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 193.595000 61.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 193.995000 61.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 194.395000 61.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.590000 194.795000 61.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 25.850000 62.110000 26.170000 ;
      LAYER met4 ;
        RECT 61.790000 25.850000 62.110000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 26.280000 62.110000 26.600000 ;
      LAYER met4 ;
        RECT 61.790000 26.280000 62.110000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 26.710000 62.110000 27.030000 ;
      LAYER met4 ;
        RECT 61.790000 26.710000 62.110000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 27.140000 62.110000 27.460000 ;
      LAYER met4 ;
        RECT 61.790000 27.140000 62.110000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 27.570000 62.110000 27.890000 ;
      LAYER met4 ;
        RECT 61.790000 27.570000 62.110000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 28.000000 62.110000 28.320000 ;
      LAYER met4 ;
        RECT 61.790000 28.000000 62.110000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 28.430000 62.110000 28.750000 ;
      LAYER met4 ;
        RECT 61.790000 28.430000 62.110000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 28.860000 62.110000 29.180000 ;
      LAYER met4 ;
        RECT 61.790000 28.860000 62.110000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 29.290000 62.110000 29.610000 ;
      LAYER met4 ;
        RECT 61.790000 29.290000 62.110000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 29.720000 62.110000 30.040000 ;
      LAYER met4 ;
        RECT 61.790000 29.720000 62.110000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 30.150000 62.110000 30.470000 ;
      LAYER met4 ;
        RECT 61.790000 30.150000 62.110000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 195.140000 62.250000 195.460000 ;
      LAYER met4 ;
        RECT 61.930000 195.140000 62.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 195.545000 62.250000 195.865000 ;
      LAYER met4 ;
        RECT 61.930000 195.545000 62.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 195.950000 62.250000 196.270000 ;
      LAYER met4 ;
        RECT 61.930000 195.950000 62.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 196.355000 62.250000 196.675000 ;
      LAYER met4 ;
        RECT 61.930000 196.355000 62.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 196.760000 62.250000 197.080000 ;
      LAYER met4 ;
        RECT 61.930000 196.760000 62.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 197.165000 62.250000 197.485000 ;
      LAYER met4 ;
        RECT 61.930000 197.165000 62.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 197.570000 62.250000 197.890000 ;
      LAYER met4 ;
        RECT 61.930000 197.570000 62.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 197.975000 62.250000 198.295000 ;
      LAYER met4 ;
        RECT 61.930000 197.975000 62.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 198.380000 62.250000 198.700000 ;
      LAYER met4 ;
        RECT 61.930000 198.380000 62.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 198.785000 62.250000 199.105000 ;
      LAYER met4 ;
        RECT 61.930000 198.785000 62.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 199.190000 62.250000 199.510000 ;
      LAYER met4 ;
        RECT 61.930000 199.190000 62.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930000 199.595000 62.250000 199.915000 ;
      LAYER met4 ;
        RECT 61.930000 199.595000 62.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 175.995000 62.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 176.395000 62.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 176.795000 62.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 177.195000 62.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 177.595000 62.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 177.995000 62.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 178.395000 62.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 178.795000 62.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 179.195000 62.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 179.595000 62.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 179.995000 62.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 180.395000 62.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 180.795000 62.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 181.195000 62.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 181.595000 62.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 181.995000 62.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 182.395000 62.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 182.795000 62.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 183.195000 62.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 183.595000 62.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 183.995000 62.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 184.395000 62.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 184.795000 62.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 185.195000 62.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 185.595000 62.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 185.995000 62.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 186.395000 62.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 186.795000 62.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 187.195000 62.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 187.595000 62.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 187.995000 62.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 188.395000 62.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 188.795000 62.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 189.195000 62.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 189.595000 62.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 189.995000 62.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 190.395000 62.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 190.795000 62.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 191.195000 62.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 191.595000 62.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 191.995000 62.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 192.395000 62.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 192.795000 62.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 193.195000 62.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 193.595000 62.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 193.995000 62.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 194.395000 62.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.990000 194.795000 62.190000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 25.850000 62.515000 26.170000 ;
      LAYER met4 ;
        RECT 62.195000 25.850000 62.515000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 26.280000 62.515000 26.600000 ;
      LAYER met4 ;
        RECT 62.195000 26.280000 62.515000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 26.710000 62.515000 27.030000 ;
      LAYER met4 ;
        RECT 62.195000 26.710000 62.515000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 27.140000 62.515000 27.460000 ;
      LAYER met4 ;
        RECT 62.195000 27.140000 62.515000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 27.570000 62.515000 27.890000 ;
      LAYER met4 ;
        RECT 62.195000 27.570000 62.515000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 28.000000 62.515000 28.320000 ;
      LAYER met4 ;
        RECT 62.195000 28.000000 62.515000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 28.430000 62.515000 28.750000 ;
      LAYER met4 ;
        RECT 62.195000 28.430000 62.515000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 28.860000 62.515000 29.180000 ;
      LAYER met4 ;
        RECT 62.195000 28.860000 62.515000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 29.290000 62.515000 29.610000 ;
      LAYER met4 ;
        RECT 62.195000 29.290000 62.515000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 29.720000 62.515000 30.040000 ;
      LAYER met4 ;
        RECT 62.195000 29.720000 62.515000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 30.150000 62.515000 30.470000 ;
      LAYER met4 ;
        RECT 62.195000 30.150000 62.515000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 195.140000 62.650000 195.460000 ;
      LAYER met4 ;
        RECT 62.330000 195.140000 62.650000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 195.545000 62.650000 195.865000 ;
      LAYER met4 ;
        RECT 62.330000 195.545000 62.650000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 195.950000 62.650000 196.270000 ;
      LAYER met4 ;
        RECT 62.330000 195.950000 62.650000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 196.355000 62.650000 196.675000 ;
      LAYER met4 ;
        RECT 62.330000 196.355000 62.650000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 196.760000 62.650000 197.080000 ;
      LAYER met4 ;
        RECT 62.330000 196.760000 62.650000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 197.165000 62.650000 197.485000 ;
      LAYER met4 ;
        RECT 62.330000 197.165000 62.650000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 197.570000 62.650000 197.890000 ;
      LAYER met4 ;
        RECT 62.330000 197.570000 62.650000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 197.975000 62.650000 198.295000 ;
      LAYER met4 ;
        RECT 62.330000 197.975000 62.650000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 198.380000 62.650000 198.700000 ;
      LAYER met4 ;
        RECT 62.330000 198.380000 62.650000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 198.785000 62.650000 199.105000 ;
      LAYER met4 ;
        RECT 62.330000 198.785000 62.650000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 199.190000 62.650000 199.510000 ;
      LAYER met4 ;
        RECT 62.330000 199.190000 62.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330000 199.595000 62.650000 199.915000 ;
      LAYER met4 ;
        RECT 62.330000 199.595000 62.650000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 175.995000 62.590000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 176.395000 62.590000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 176.795000 62.590000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 177.195000 62.590000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 177.595000 62.590000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 177.995000 62.590000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 178.395000 62.590000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 178.795000 62.590000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 179.195000 62.590000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 179.595000 62.590000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 179.995000 62.590000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 180.395000 62.590000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 180.795000 62.590000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 181.195000 62.590000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 181.595000 62.590000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 181.995000 62.590000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 182.395000 62.590000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 182.795000 62.590000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 183.195000 62.590000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 183.595000 62.590000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 183.995000 62.590000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 184.395000 62.590000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 184.795000 62.590000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 185.195000 62.590000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 185.595000 62.590000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 185.995000 62.590000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 186.395000 62.590000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 186.795000 62.590000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 187.195000 62.590000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 187.595000 62.590000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 187.995000 62.590000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 188.395000 62.590000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 188.795000 62.590000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 189.195000 62.590000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 189.595000 62.590000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 189.995000 62.590000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 190.395000 62.590000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 190.795000 62.590000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 191.195000 62.590000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 191.595000 62.590000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 191.995000 62.590000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 192.395000 62.590000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 192.795000 62.590000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 193.195000 62.590000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 193.595000 62.590000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 193.995000 62.590000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 194.395000 62.590000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.390000 194.795000 62.590000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 25.850000 62.920000 26.170000 ;
      LAYER met4 ;
        RECT 62.600000 25.850000 62.920000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 26.280000 62.920000 26.600000 ;
      LAYER met4 ;
        RECT 62.600000 26.280000 62.920000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 26.710000 62.920000 27.030000 ;
      LAYER met4 ;
        RECT 62.600000 26.710000 62.920000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 27.140000 62.920000 27.460000 ;
      LAYER met4 ;
        RECT 62.600000 27.140000 62.920000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 27.570000 62.920000 27.890000 ;
      LAYER met4 ;
        RECT 62.600000 27.570000 62.920000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 28.000000 62.920000 28.320000 ;
      LAYER met4 ;
        RECT 62.600000 28.000000 62.920000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 28.430000 62.920000 28.750000 ;
      LAYER met4 ;
        RECT 62.600000 28.430000 62.920000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 28.860000 62.920000 29.180000 ;
      LAYER met4 ;
        RECT 62.600000 28.860000 62.920000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 29.290000 62.920000 29.610000 ;
      LAYER met4 ;
        RECT 62.600000 29.290000 62.920000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 29.720000 62.920000 30.040000 ;
      LAYER met4 ;
        RECT 62.600000 29.720000 62.920000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 30.150000 62.920000 30.470000 ;
      LAYER met4 ;
        RECT 62.600000 30.150000 62.920000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 195.140000 63.050000 195.460000 ;
      LAYER met4 ;
        RECT 62.730000 195.140000 63.050000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 195.545000 63.050000 195.865000 ;
      LAYER met4 ;
        RECT 62.730000 195.545000 63.050000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 195.950000 63.050000 196.270000 ;
      LAYER met4 ;
        RECT 62.730000 195.950000 63.050000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 196.355000 63.050000 196.675000 ;
      LAYER met4 ;
        RECT 62.730000 196.355000 63.050000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 196.760000 63.050000 197.080000 ;
      LAYER met4 ;
        RECT 62.730000 196.760000 63.050000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 197.165000 63.050000 197.485000 ;
      LAYER met4 ;
        RECT 62.730000 197.165000 63.050000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 197.570000 63.050000 197.890000 ;
      LAYER met4 ;
        RECT 62.730000 197.570000 63.050000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 197.975000 63.050000 198.295000 ;
      LAYER met4 ;
        RECT 62.730000 197.975000 63.050000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 198.380000 63.050000 198.700000 ;
      LAYER met4 ;
        RECT 62.730000 198.380000 63.050000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 198.785000 63.050000 199.105000 ;
      LAYER met4 ;
        RECT 62.730000 198.785000 63.050000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 199.190000 63.050000 199.510000 ;
      LAYER met4 ;
        RECT 62.730000 199.190000 63.050000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730000 199.595000 63.050000 199.915000 ;
      LAYER met4 ;
        RECT 62.730000 199.595000 63.050000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 175.995000 62.990000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 176.395000 62.990000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 176.795000 62.990000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 177.195000 62.990000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 177.595000 62.990000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 177.995000 62.990000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 178.395000 62.990000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 178.795000 62.990000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 179.195000 62.990000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 179.595000 62.990000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 179.995000 62.990000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 180.395000 62.990000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 180.795000 62.990000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 181.195000 62.990000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 181.595000 62.990000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 181.995000 62.990000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 182.395000 62.990000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 182.795000 62.990000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 183.195000 62.990000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 183.595000 62.990000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 183.995000 62.990000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 184.395000 62.990000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 184.795000 62.990000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 185.195000 62.990000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 185.595000 62.990000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 185.995000 62.990000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 186.395000 62.990000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 186.795000 62.990000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 187.195000 62.990000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 187.595000 62.990000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 187.995000 62.990000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 188.395000 62.990000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 188.795000 62.990000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 189.195000 62.990000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 189.595000 62.990000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 189.995000 62.990000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 190.395000 62.990000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 190.795000 62.990000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 191.195000 62.990000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 191.595000 62.990000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 191.995000 62.990000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 192.395000 62.990000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 192.795000 62.990000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 193.195000 62.990000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 193.595000 62.990000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 193.995000 62.990000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 194.395000 62.990000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.790000 194.795000 62.990000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 25.850000 63.325000 26.170000 ;
      LAYER met4 ;
        RECT 63.005000 25.850000 63.325000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 26.280000 63.325000 26.600000 ;
      LAYER met4 ;
        RECT 63.005000 26.280000 63.325000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 26.710000 63.325000 27.030000 ;
      LAYER met4 ;
        RECT 63.005000 26.710000 63.325000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 27.140000 63.325000 27.460000 ;
      LAYER met4 ;
        RECT 63.005000 27.140000 63.325000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 27.570000 63.325000 27.890000 ;
      LAYER met4 ;
        RECT 63.005000 27.570000 63.325000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 28.000000 63.325000 28.320000 ;
      LAYER met4 ;
        RECT 63.005000 28.000000 63.325000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 28.430000 63.325000 28.750000 ;
      LAYER met4 ;
        RECT 63.005000 28.430000 63.325000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 28.860000 63.325000 29.180000 ;
      LAYER met4 ;
        RECT 63.005000 28.860000 63.325000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 29.290000 63.325000 29.610000 ;
      LAYER met4 ;
        RECT 63.005000 29.290000 63.325000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 29.720000 63.325000 30.040000 ;
      LAYER met4 ;
        RECT 63.005000 29.720000 63.325000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 30.150000 63.325000 30.470000 ;
      LAYER met4 ;
        RECT 63.005000 30.150000 63.325000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 195.140000 63.450000 195.460000 ;
      LAYER met4 ;
        RECT 63.130000 195.140000 63.450000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 195.545000 63.450000 195.865000 ;
      LAYER met4 ;
        RECT 63.130000 195.545000 63.450000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 195.950000 63.450000 196.270000 ;
      LAYER met4 ;
        RECT 63.130000 195.950000 63.450000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 196.355000 63.450000 196.675000 ;
      LAYER met4 ;
        RECT 63.130000 196.355000 63.450000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 196.760000 63.450000 197.080000 ;
      LAYER met4 ;
        RECT 63.130000 196.760000 63.450000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 197.165000 63.450000 197.485000 ;
      LAYER met4 ;
        RECT 63.130000 197.165000 63.450000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 197.570000 63.450000 197.890000 ;
      LAYER met4 ;
        RECT 63.130000 197.570000 63.450000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 197.975000 63.450000 198.295000 ;
      LAYER met4 ;
        RECT 63.130000 197.975000 63.450000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 198.380000 63.450000 198.700000 ;
      LAYER met4 ;
        RECT 63.130000 198.380000 63.450000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 198.785000 63.450000 199.105000 ;
      LAYER met4 ;
        RECT 63.130000 198.785000 63.450000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 199.190000 63.450000 199.510000 ;
      LAYER met4 ;
        RECT 63.130000 199.190000 63.450000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130000 199.595000 63.450000 199.915000 ;
      LAYER met4 ;
        RECT 63.130000 199.595000 63.450000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 175.995000 63.390000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 176.395000 63.390000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 176.795000 63.390000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 177.195000 63.390000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 177.595000 63.390000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 177.995000 63.390000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 178.395000 63.390000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 178.795000 63.390000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 179.195000 63.390000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 179.595000 63.390000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 179.995000 63.390000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 180.395000 63.390000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 180.795000 63.390000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 181.195000 63.390000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 181.595000 63.390000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 181.995000 63.390000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 182.395000 63.390000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 182.795000 63.390000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 183.195000 63.390000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 183.595000 63.390000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 183.995000 63.390000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 184.395000 63.390000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 184.795000 63.390000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 185.195000 63.390000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 185.595000 63.390000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 185.995000 63.390000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 186.395000 63.390000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 186.795000 63.390000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 187.195000 63.390000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 187.595000 63.390000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 187.995000 63.390000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 188.395000 63.390000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 188.795000 63.390000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 189.195000 63.390000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 189.595000 63.390000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 189.995000 63.390000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 190.395000 63.390000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 190.795000 63.390000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 191.195000 63.390000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 191.595000 63.390000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 191.995000 63.390000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 192.395000 63.390000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 192.795000 63.390000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 193.195000 63.390000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 193.595000 63.390000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 193.995000 63.390000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 194.395000 63.390000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 194.795000 63.390000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 25.850000 63.730000 26.170000 ;
      LAYER met4 ;
        RECT 63.410000 25.850000 63.730000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 26.280000 63.730000 26.600000 ;
      LAYER met4 ;
        RECT 63.410000 26.280000 63.730000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 26.710000 63.730000 27.030000 ;
      LAYER met4 ;
        RECT 63.410000 26.710000 63.730000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 27.140000 63.730000 27.460000 ;
      LAYER met4 ;
        RECT 63.410000 27.140000 63.730000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 27.570000 63.730000 27.890000 ;
      LAYER met4 ;
        RECT 63.410000 27.570000 63.730000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 28.000000 63.730000 28.320000 ;
      LAYER met4 ;
        RECT 63.410000 28.000000 63.730000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 28.430000 63.730000 28.750000 ;
      LAYER met4 ;
        RECT 63.410000 28.430000 63.730000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 28.860000 63.730000 29.180000 ;
      LAYER met4 ;
        RECT 63.410000 28.860000 63.730000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 29.290000 63.730000 29.610000 ;
      LAYER met4 ;
        RECT 63.410000 29.290000 63.730000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 29.720000 63.730000 30.040000 ;
      LAYER met4 ;
        RECT 63.410000 29.720000 63.730000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 30.150000 63.730000 30.470000 ;
      LAYER met4 ;
        RECT 63.410000 30.150000 63.730000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 195.140000 63.850000 195.460000 ;
      LAYER met4 ;
        RECT 63.530000 195.140000 63.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 195.545000 63.850000 195.865000 ;
      LAYER met4 ;
        RECT 63.530000 195.545000 63.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 195.950000 63.850000 196.270000 ;
      LAYER met4 ;
        RECT 63.530000 195.950000 63.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 196.355000 63.850000 196.675000 ;
      LAYER met4 ;
        RECT 63.530000 196.355000 63.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 196.760000 63.850000 197.080000 ;
      LAYER met4 ;
        RECT 63.530000 196.760000 63.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 197.165000 63.850000 197.485000 ;
      LAYER met4 ;
        RECT 63.530000 197.165000 63.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 197.570000 63.850000 197.890000 ;
      LAYER met4 ;
        RECT 63.530000 197.570000 63.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 197.975000 63.850000 198.295000 ;
      LAYER met4 ;
        RECT 63.530000 197.975000 63.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 198.380000 63.850000 198.700000 ;
      LAYER met4 ;
        RECT 63.530000 198.380000 63.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 198.785000 63.850000 199.105000 ;
      LAYER met4 ;
        RECT 63.530000 198.785000 63.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 199.190000 63.850000 199.510000 ;
      LAYER met4 ;
        RECT 63.530000 199.190000 63.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530000 199.595000 63.850000 199.915000 ;
      LAYER met4 ;
        RECT 63.530000 199.595000 63.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 175.995000 63.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 176.395000 63.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 176.795000 63.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 177.195000 63.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 177.595000 63.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 177.995000 63.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 178.395000 63.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 178.795000 63.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 179.195000 63.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 179.595000 63.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 179.995000 63.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 180.395000 63.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 180.795000 63.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 181.195000 63.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 181.595000 63.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 181.995000 63.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 182.395000 63.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 182.795000 63.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 183.195000 63.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 183.595000 63.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 183.995000 63.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 184.395000 63.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 184.795000 63.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 185.195000 63.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 185.595000 63.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 185.995000 63.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 186.395000 63.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 186.795000 63.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 187.195000 63.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 187.595000 63.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 187.995000 63.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 188.395000 63.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 188.795000 63.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 189.195000 63.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 189.595000 63.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 189.995000 63.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 190.395000 63.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 190.795000 63.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 191.195000 63.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 191.595000 63.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 191.995000 63.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 192.395000 63.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 192.795000 63.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 193.195000 63.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 193.595000 63.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 193.995000 63.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 194.395000 63.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.590000 194.795000 63.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 25.850000 64.135000 26.170000 ;
      LAYER met4 ;
        RECT 63.815000 25.850000 64.135000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 26.280000 64.135000 26.600000 ;
      LAYER met4 ;
        RECT 63.815000 26.280000 64.135000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 26.710000 64.135000 27.030000 ;
      LAYER met4 ;
        RECT 63.815000 26.710000 64.135000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 27.140000 64.135000 27.460000 ;
      LAYER met4 ;
        RECT 63.815000 27.140000 64.135000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 27.570000 64.135000 27.890000 ;
      LAYER met4 ;
        RECT 63.815000 27.570000 64.135000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 28.000000 64.135000 28.320000 ;
      LAYER met4 ;
        RECT 63.815000 28.000000 64.135000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 28.430000 64.135000 28.750000 ;
      LAYER met4 ;
        RECT 63.815000 28.430000 64.135000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 28.860000 64.135000 29.180000 ;
      LAYER met4 ;
        RECT 63.815000 28.860000 64.135000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 29.290000 64.135000 29.610000 ;
      LAYER met4 ;
        RECT 63.815000 29.290000 64.135000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 29.720000 64.135000 30.040000 ;
      LAYER met4 ;
        RECT 63.815000 29.720000 64.135000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 30.150000 64.135000 30.470000 ;
      LAYER met4 ;
        RECT 63.815000 30.150000 64.135000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 195.140000 64.250000 195.460000 ;
      LAYER met4 ;
        RECT 63.930000 195.140000 64.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 195.545000 64.250000 195.865000 ;
      LAYER met4 ;
        RECT 63.930000 195.545000 64.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 195.950000 64.250000 196.270000 ;
      LAYER met4 ;
        RECT 63.930000 195.950000 64.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 196.355000 64.250000 196.675000 ;
      LAYER met4 ;
        RECT 63.930000 196.355000 64.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 196.760000 64.250000 197.080000 ;
      LAYER met4 ;
        RECT 63.930000 196.760000 64.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 197.165000 64.250000 197.485000 ;
      LAYER met4 ;
        RECT 63.930000 197.165000 64.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 197.570000 64.250000 197.890000 ;
      LAYER met4 ;
        RECT 63.930000 197.570000 64.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 197.975000 64.250000 198.295000 ;
      LAYER met4 ;
        RECT 63.930000 197.975000 64.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 198.380000 64.250000 198.700000 ;
      LAYER met4 ;
        RECT 63.930000 198.380000 64.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 198.785000 64.250000 199.105000 ;
      LAYER met4 ;
        RECT 63.930000 198.785000 64.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 199.190000 64.250000 199.510000 ;
      LAYER met4 ;
        RECT 63.930000 199.190000 64.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930000 199.595000 64.250000 199.915000 ;
      LAYER met4 ;
        RECT 63.930000 199.595000 64.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 175.995000 64.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 176.395000 64.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 176.795000 64.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 177.195000 64.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 177.595000 64.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 177.995000 64.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 178.395000 64.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 178.795000 64.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 179.195000 64.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 179.595000 64.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 179.995000 64.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 180.395000 64.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 180.795000 64.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 181.195000 64.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 181.595000 64.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 181.995000 64.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 182.395000 64.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 182.795000 64.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 183.195000 64.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 183.595000 64.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 183.995000 64.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 184.395000 64.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 184.795000 64.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 185.195000 64.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 185.595000 64.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 185.995000 64.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 186.395000 64.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 186.795000 64.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 187.195000 64.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 187.595000 64.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 187.995000 64.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 188.395000 64.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 188.795000 64.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 189.195000 64.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 189.595000 64.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 189.995000 64.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 190.395000 64.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 190.795000 64.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 191.195000 64.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 191.595000 64.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 191.995000 64.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 192.395000 64.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 192.795000 64.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 193.195000 64.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 193.595000 64.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 193.995000 64.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 194.395000 64.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.990000 194.795000 64.190000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 25.850000 64.540000 26.170000 ;
      LAYER met4 ;
        RECT 64.220000 25.850000 64.540000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 26.280000 64.540000 26.600000 ;
      LAYER met4 ;
        RECT 64.220000 26.280000 64.540000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 26.710000 64.540000 27.030000 ;
      LAYER met4 ;
        RECT 64.220000 26.710000 64.540000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 27.140000 64.540000 27.460000 ;
      LAYER met4 ;
        RECT 64.220000 27.140000 64.540000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 27.570000 64.540000 27.890000 ;
      LAYER met4 ;
        RECT 64.220000 27.570000 64.540000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 28.000000 64.540000 28.320000 ;
      LAYER met4 ;
        RECT 64.220000 28.000000 64.540000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 28.430000 64.540000 28.750000 ;
      LAYER met4 ;
        RECT 64.220000 28.430000 64.540000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 28.860000 64.540000 29.180000 ;
      LAYER met4 ;
        RECT 64.220000 28.860000 64.540000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 29.290000 64.540000 29.610000 ;
      LAYER met4 ;
        RECT 64.220000 29.290000 64.540000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 29.720000 64.540000 30.040000 ;
      LAYER met4 ;
        RECT 64.220000 29.720000 64.540000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 30.150000 64.540000 30.470000 ;
      LAYER met4 ;
        RECT 64.220000 30.150000 64.540000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 195.140000 64.650000 195.460000 ;
      LAYER met4 ;
        RECT 64.330000 195.140000 64.650000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 195.545000 64.650000 195.865000 ;
      LAYER met4 ;
        RECT 64.330000 195.545000 64.650000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 195.950000 64.650000 196.270000 ;
      LAYER met4 ;
        RECT 64.330000 195.950000 64.650000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 196.355000 64.650000 196.675000 ;
      LAYER met4 ;
        RECT 64.330000 196.355000 64.650000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 196.760000 64.650000 197.080000 ;
      LAYER met4 ;
        RECT 64.330000 196.760000 64.650000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 197.165000 64.650000 197.485000 ;
      LAYER met4 ;
        RECT 64.330000 197.165000 64.650000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 197.570000 64.650000 197.890000 ;
      LAYER met4 ;
        RECT 64.330000 197.570000 64.650000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 197.975000 64.650000 198.295000 ;
      LAYER met4 ;
        RECT 64.330000 197.975000 64.650000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 198.380000 64.650000 198.700000 ;
      LAYER met4 ;
        RECT 64.330000 198.380000 64.650000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 198.785000 64.650000 199.105000 ;
      LAYER met4 ;
        RECT 64.330000 198.785000 64.650000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 199.190000 64.650000 199.510000 ;
      LAYER met4 ;
        RECT 64.330000 199.190000 64.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330000 199.595000 64.650000 199.915000 ;
      LAYER met4 ;
        RECT 64.330000 199.595000 64.650000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 175.995000 64.590000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 176.395000 64.590000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 176.795000 64.590000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 177.195000 64.590000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 177.595000 64.590000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 177.995000 64.590000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 178.395000 64.590000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 178.795000 64.590000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 179.195000 64.590000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 179.595000 64.590000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 179.995000 64.590000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 180.395000 64.590000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 180.795000 64.590000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 181.195000 64.590000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 181.595000 64.590000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 181.995000 64.590000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 182.395000 64.590000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 182.795000 64.590000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 183.195000 64.590000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 183.595000 64.590000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 183.995000 64.590000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 184.395000 64.590000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 184.795000 64.590000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 185.195000 64.590000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 185.595000 64.590000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 185.995000 64.590000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 186.395000 64.590000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 186.795000 64.590000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 187.195000 64.590000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 187.595000 64.590000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 187.995000 64.590000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 188.395000 64.590000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 188.795000 64.590000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 189.195000 64.590000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 189.595000 64.590000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 189.995000 64.590000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 190.395000 64.590000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 190.795000 64.590000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 191.195000 64.590000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 191.595000 64.590000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 191.995000 64.590000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 192.395000 64.590000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 192.795000 64.590000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 193.195000 64.590000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 193.595000 64.590000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 193.995000 64.590000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 194.395000 64.590000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.390000 194.795000 64.590000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 25.850000 64.945000 26.170000 ;
      LAYER met4 ;
        RECT 64.625000 25.850000 64.945000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 26.280000 64.945000 26.600000 ;
      LAYER met4 ;
        RECT 64.625000 26.280000 64.945000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 26.710000 64.945000 27.030000 ;
      LAYER met4 ;
        RECT 64.625000 26.710000 64.945000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 27.140000 64.945000 27.460000 ;
      LAYER met4 ;
        RECT 64.625000 27.140000 64.945000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 27.570000 64.945000 27.890000 ;
      LAYER met4 ;
        RECT 64.625000 27.570000 64.945000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 28.000000 64.945000 28.320000 ;
      LAYER met4 ;
        RECT 64.625000 28.000000 64.945000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 28.430000 64.945000 28.750000 ;
      LAYER met4 ;
        RECT 64.625000 28.430000 64.945000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 28.860000 64.945000 29.180000 ;
      LAYER met4 ;
        RECT 64.625000 28.860000 64.945000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 29.290000 64.945000 29.610000 ;
      LAYER met4 ;
        RECT 64.625000 29.290000 64.945000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 29.720000 64.945000 30.040000 ;
      LAYER met4 ;
        RECT 64.625000 29.720000 64.945000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 30.150000 64.945000 30.470000 ;
      LAYER met4 ;
        RECT 64.625000 30.150000 64.945000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 195.140000 65.050000 195.460000 ;
      LAYER met4 ;
        RECT 64.730000 195.140000 65.050000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 195.545000 65.050000 195.865000 ;
      LAYER met4 ;
        RECT 64.730000 195.545000 65.050000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 195.950000 65.050000 196.270000 ;
      LAYER met4 ;
        RECT 64.730000 195.950000 65.050000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 196.355000 65.050000 196.675000 ;
      LAYER met4 ;
        RECT 64.730000 196.355000 65.050000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 196.760000 65.050000 197.080000 ;
      LAYER met4 ;
        RECT 64.730000 196.760000 65.050000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 197.165000 65.050000 197.485000 ;
      LAYER met4 ;
        RECT 64.730000 197.165000 65.050000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 197.570000 65.050000 197.890000 ;
      LAYER met4 ;
        RECT 64.730000 197.570000 65.050000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 197.975000 65.050000 198.295000 ;
      LAYER met4 ;
        RECT 64.730000 197.975000 65.050000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 198.380000 65.050000 198.700000 ;
      LAYER met4 ;
        RECT 64.730000 198.380000 65.050000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 198.785000 65.050000 199.105000 ;
      LAYER met4 ;
        RECT 64.730000 198.785000 65.050000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 199.190000 65.050000 199.510000 ;
      LAYER met4 ;
        RECT 64.730000 199.190000 65.050000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730000 199.595000 65.050000 199.915000 ;
      LAYER met4 ;
        RECT 64.730000 199.595000 65.050000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 175.995000 64.990000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 176.395000 64.990000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 176.795000 64.990000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 177.195000 64.990000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 177.595000 64.990000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 177.995000 64.990000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 178.395000 64.990000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 178.795000 64.990000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 179.195000 64.990000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 179.595000 64.990000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 179.995000 64.990000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 180.395000 64.990000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 180.795000 64.990000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 181.195000 64.990000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 181.595000 64.990000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 181.995000 64.990000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 182.395000 64.990000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 182.795000 64.990000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 183.195000 64.990000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 183.595000 64.990000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 183.995000 64.990000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 184.395000 64.990000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 184.795000 64.990000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 185.195000 64.990000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 185.595000 64.990000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 185.995000 64.990000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 186.395000 64.990000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 186.795000 64.990000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 187.195000 64.990000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 187.595000 64.990000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 187.995000 64.990000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 188.395000 64.990000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 188.795000 64.990000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 189.195000 64.990000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 189.595000 64.990000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 189.995000 64.990000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 190.395000 64.990000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 190.795000 64.990000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 191.195000 64.990000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 191.595000 64.990000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 191.995000 64.990000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 192.395000 64.990000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 192.795000 64.990000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 193.195000 64.990000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 193.595000 64.990000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 193.995000 64.990000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 194.395000 64.990000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.790000 194.795000 64.990000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 25.850000 65.350000 26.170000 ;
      LAYER met4 ;
        RECT 65.030000 25.850000 65.350000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 26.280000 65.350000 26.600000 ;
      LAYER met4 ;
        RECT 65.030000 26.280000 65.350000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 26.710000 65.350000 27.030000 ;
      LAYER met4 ;
        RECT 65.030000 26.710000 65.350000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 27.140000 65.350000 27.460000 ;
      LAYER met4 ;
        RECT 65.030000 27.140000 65.350000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 27.570000 65.350000 27.890000 ;
      LAYER met4 ;
        RECT 65.030000 27.570000 65.350000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 28.000000 65.350000 28.320000 ;
      LAYER met4 ;
        RECT 65.030000 28.000000 65.350000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 28.430000 65.350000 28.750000 ;
      LAYER met4 ;
        RECT 65.030000 28.430000 65.350000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 28.860000 65.350000 29.180000 ;
      LAYER met4 ;
        RECT 65.030000 28.860000 65.350000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 29.290000 65.350000 29.610000 ;
      LAYER met4 ;
        RECT 65.030000 29.290000 65.350000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 29.720000 65.350000 30.040000 ;
      LAYER met4 ;
        RECT 65.030000 29.720000 65.350000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 30.150000 65.350000 30.470000 ;
      LAYER met4 ;
        RECT 65.030000 30.150000 65.350000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 195.140000 65.450000 195.460000 ;
      LAYER met4 ;
        RECT 65.130000 195.140000 65.450000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 195.545000 65.450000 195.865000 ;
      LAYER met4 ;
        RECT 65.130000 195.545000 65.450000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 195.950000 65.450000 196.270000 ;
      LAYER met4 ;
        RECT 65.130000 195.950000 65.450000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 196.355000 65.450000 196.675000 ;
      LAYER met4 ;
        RECT 65.130000 196.355000 65.450000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 196.760000 65.450000 197.080000 ;
      LAYER met4 ;
        RECT 65.130000 196.760000 65.450000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 197.165000 65.450000 197.485000 ;
      LAYER met4 ;
        RECT 65.130000 197.165000 65.450000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 197.570000 65.450000 197.890000 ;
      LAYER met4 ;
        RECT 65.130000 197.570000 65.450000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 197.975000 65.450000 198.295000 ;
      LAYER met4 ;
        RECT 65.130000 197.975000 65.450000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 198.380000 65.450000 198.700000 ;
      LAYER met4 ;
        RECT 65.130000 198.380000 65.450000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 198.785000 65.450000 199.105000 ;
      LAYER met4 ;
        RECT 65.130000 198.785000 65.450000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 199.190000 65.450000 199.510000 ;
      LAYER met4 ;
        RECT 65.130000 199.190000 65.450000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130000 199.595000 65.450000 199.915000 ;
      LAYER met4 ;
        RECT 65.130000 199.595000 65.450000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 175.995000 65.390000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 176.395000 65.390000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 176.795000 65.390000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 177.195000 65.390000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 177.595000 65.390000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 177.995000 65.390000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 178.395000 65.390000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 178.795000 65.390000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 179.195000 65.390000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 179.595000 65.390000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 179.995000 65.390000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 180.395000 65.390000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 180.795000 65.390000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 181.195000 65.390000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 181.595000 65.390000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 181.995000 65.390000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 182.395000 65.390000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 182.795000 65.390000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 183.195000 65.390000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 183.595000 65.390000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 183.995000 65.390000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 184.395000 65.390000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 184.795000 65.390000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 185.195000 65.390000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 185.595000 65.390000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 185.995000 65.390000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 186.395000 65.390000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 186.795000 65.390000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 187.195000 65.390000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 187.595000 65.390000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 187.995000 65.390000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 188.395000 65.390000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 188.795000 65.390000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 189.195000 65.390000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 189.595000 65.390000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 189.995000 65.390000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 190.395000 65.390000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 190.795000 65.390000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 191.195000 65.390000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 191.595000 65.390000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 191.995000 65.390000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 192.395000 65.390000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 192.795000 65.390000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 193.195000 65.390000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 193.595000 65.390000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 193.995000 65.390000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 194.395000 65.390000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.190000 194.795000 65.390000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 25.850000 65.755000 26.170000 ;
      LAYER met4 ;
        RECT 65.435000 25.850000 65.755000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 26.280000 65.755000 26.600000 ;
      LAYER met4 ;
        RECT 65.435000 26.280000 65.755000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 26.710000 65.755000 27.030000 ;
      LAYER met4 ;
        RECT 65.435000 26.710000 65.755000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 27.140000 65.755000 27.460000 ;
      LAYER met4 ;
        RECT 65.435000 27.140000 65.755000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 27.570000 65.755000 27.890000 ;
      LAYER met4 ;
        RECT 65.435000 27.570000 65.755000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 28.000000 65.755000 28.320000 ;
      LAYER met4 ;
        RECT 65.435000 28.000000 65.755000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 28.430000 65.755000 28.750000 ;
      LAYER met4 ;
        RECT 65.435000 28.430000 65.755000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 28.860000 65.755000 29.180000 ;
      LAYER met4 ;
        RECT 65.435000 28.860000 65.755000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 29.290000 65.755000 29.610000 ;
      LAYER met4 ;
        RECT 65.435000 29.290000 65.755000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 29.720000 65.755000 30.040000 ;
      LAYER met4 ;
        RECT 65.435000 29.720000 65.755000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 30.150000 65.755000 30.470000 ;
      LAYER met4 ;
        RECT 65.435000 30.150000 65.755000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 195.140000 65.850000 195.460000 ;
      LAYER met4 ;
        RECT 65.530000 195.140000 65.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 195.545000 65.850000 195.865000 ;
      LAYER met4 ;
        RECT 65.530000 195.545000 65.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 195.950000 65.850000 196.270000 ;
      LAYER met4 ;
        RECT 65.530000 195.950000 65.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 196.355000 65.850000 196.675000 ;
      LAYER met4 ;
        RECT 65.530000 196.355000 65.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 196.760000 65.850000 197.080000 ;
      LAYER met4 ;
        RECT 65.530000 196.760000 65.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 197.165000 65.850000 197.485000 ;
      LAYER met4 ;
        RECT 65.530000 197.165000 65.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 197.570000 65.850000 197.890000 ;
      LAYER met4 ;
        RECT 65.530000 197.570000 65.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 197.975000 65.850000 198.295000 ;
      LAYER met4 ;
        RECT 65.530000 197.975000 65.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 198.380000 65.850000 198.700000 ;
      LAYER met4 ;
        RECT 65.530000 198.380000 65.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 198.785000 65.850000 199.105000 ;
      LAYER met4 ;
        RECT 65.530000 198.785000 65.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 199.190000 65.850000 199.510000 ;
      LAYER met4 ;
        RECT 65.530000 199.190000 65.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530000 199.595000 65.850000 199.915000 ;
      LAYER met4 ;
        RECT 65.530000 199.595000 65.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 175.995000 65.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 176.395000 65.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 176.795000 65.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 177.195000 65.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 177.595000 65.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 177.995000 65.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 178.395000 65.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 178.795000 65.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 179.195000 65.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 179.595000 65.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 179.995000 65.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 180.395000 65.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 180.795000 65.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 181.195000 65.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 181.595000 65.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 181.995000 65.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 182.395000 65.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 182.795000 65.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 183.195000 65.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 183.595000 65.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 183.995000 65.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 184.395000 65.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 184.795000 65.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 185.195000 65.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 185.595000 65.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 185.995000 65.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 186.395000 65.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 186.795000 65.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 187.195000 65.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 187.595000 65.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 187.995000 65.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 188.395000 65.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 188.795000 65.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 189.195000 65.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 189.595000 65.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 189.995000 65.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 190.395000 65.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 190.795000 65.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 191.195000 65.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 191.595000 65.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 191.995000 65.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 192.395000 65.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 192.795000 65.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 193.195000 65.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 193.595000 65.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 193.995000 65.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 194.395000 65.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 194.795000 65.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 25.850000 66.160000 26.170000 ;
      LAYER met4 ;
        RECT 65.840000 25.850000 66.160000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 26.280000 66.160000 26.600000 ;
      LAYER met4 ;
        RECT 65.840000 26.280000 66.160000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 26.710000 66.160000 27.030000 ;
      LAYER met4 ;
        RECT 65.840000 26.710000 66.160000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 27.140000 66.160000 27.460000 ;
      LAYER met4 ;
        RECT 65.840000 27.140000 66.160000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 27.570000 66.160000 27.890000 ;
      LAYER met4 ;
        RECT 65.840000 27.570000 66.160000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 28.000000 66.160000 28.320000 ;
      LAYER met4 ;
        RECT 65.840000 28.000000 66.160000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 28.430000 66.160000 28.750000 ;
      LAYER met4 ;
        RECT 65.840000 28.430000 66.160000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 28.860000 66.160000 29.180000 ;
      LAYER met4 ;
        RECT 65.840000 28.860000 66.160000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 29.290000 66.160000 29.610000 ;
      LAYER met4 ;
        RECT 65.840000 29.290000 66.160000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 29.720000 66.160000 30.040000 ;
      LAYER met4 ;
        RECT 65.840000 29.720000 66.160000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 30.150000 66.160000 30.470000 ;
      LAYER met4 ;
        RECT 65.840000 30.150000 66.160000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 195.140000 66.250000 195.460000 ;
      LAYER met4 ;
        RECT 65.930000 195.140000 66.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 195.545000 66.250000 195.865000 ;
      LAYER met4 ;
        RECT 65.930000 195.545000 66.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 195.950000 66.250000 196.270000 ;
      LAYER met4 ;
        RECT 65.930000 195.950000 66.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 196.355000 66.250000 196.675000 ;
      LAYER met4 ;
        RECT 65.930000 196.355000 66.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 196.760000 66.250000 197.080000 ;
      LAYER met4 ;
        RECT 65.930000 196.760000 66.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 197.165000 66.250000 197.485000 ;
      LAYER met4 ;
        RECT 65.930000 197.165000 66.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 197.570000 66.250000 197.890000 ;
      LAYER met4 ;
        RECT 65.930000 197.570000 66.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 197.975000 66.250000 198.295000 ;
      LAYER met4 ;
        RECT 65.930000 197.975000 66.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 198.380000 66.250000 198.700000 ;
      LAYER met4 ;
        RECT 65.930000 198.380000 66.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 198.785000 66.250000 199.105000 ;
      LAYER met4 ;
        RECT 65.930000 198.785000 66.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 199.190000 66.250000 199.510000 ;
      LAYER met4 ;
        RECT 65.930000 199.190000 66.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930000 199.595000 66.250000 199.915000 ;
      LAYER met4 ;
        RECT 65.930000 199.595000 66.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 175.995000 66.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 176.395000 66.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 176.795000 66.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 177.195000 66.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 177.595000 66.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 177.995000 66.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 178.395000 66.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 178.795000 66.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 179.195000 66.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 179.595000 66.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 179.995000 66.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 180.395000 66.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 180.795000 66.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 181.195000 66.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 181.595000 66.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 181.995000 66.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 182.395000 66.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 182.795000 66.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 183.195000 66.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 183.595000 66.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 183.995000 66.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 184.395000 66.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 184.795000 66.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 185.195000 66.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 185.595000 66.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 185.995000 66.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 186.395000 66.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 186.795000 66.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 187.195000 66.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 187.595000 66.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 187.995000 66.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 188.395000 66.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 188.795000 66.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 189.195000 66.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 189.595000 66.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 189.995000 66.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 190.395000 66.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 190.795000 66.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 191.195000 66.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 191.595000 66.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 191.995000 66.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 192.395000 66.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 192.795000 66.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 193.195000 66.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 193.595000 66.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 193.995000 66.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 194.395000 66.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 194.795000 66.190000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 25.850000 66.565000 26.170000 ;
      LAYER met4 ;
        RECT 66.245000 25.850000 66.565000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 26.280000 66.565000 26.600000 ;
      LAYER met4 ;
        RECT 66.245000 26.280000 66.565000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 26.710000 66.565000 27.030000 ;
      LAYER met4 ;
        RECT 66.245000 26.710000 66.565000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 27.140000 66.565000 27.460000 ;
      LAYER met4 ;
        RECT 66.245000 27.140000 66.565000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 27.570000 66.565000 27.890000 ;
      LAYER met4 ;
        RECT 66.245000 27.570000 66.565000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 28.000000 66.565000 28.320000 ;
      LAYER met4 ;
        RECT 66.245000 28.000000 66.565000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 28.430000 66.565000 28.750000 ;
      LAYER met4 ;
        RECT 66.245000 28.430000 66.565000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 28.860000 66.565000 29.180000 ;
      LAYER met4 ;
        RECT 66.245000 28.860000 66.565000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 29.290000 66.565000 29.610000 ;
      LAYER met4 ;
        RECT 66.245000 29.290000 66.565000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 29.720000 66.565000 30.040000 ;
      LAYER met4 ;
        RECT 66.245000 29.720000 66.565000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 30.150000 66.565000 30.470000 ;
      LAYER met4 ;
        RECT 66.245000 30.150000 66.565000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 195.140000 66.650000 195.460000 ;
      LAYER met4 ;
        RECT 66.330000 195.140000 66.650000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 195.545000 66.650000 195.865000 ;
      LAYER met4 ;
        RECT 66.330000 195.545000 66.650000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 195.950000 66.650000 196.270000 ;
      LAYER met4 ;
        RECT 66.330000 195.950000 66.650000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 196.355000 66.650000 196.675000 ;
      LAYER met4 ;
        RECT 66.330000 196.355000 66.650000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 196.760000 66.650000 197.080000 ;
      LAYER met4 ;
        RECT 66.330000 196.760000 66.650000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 197.165000 66.650000 197.485000 ;
      LAYER met4 ;
        RECT 66.330000 197.165000 66.650000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 197.570000 66.650000 197.890000 ;
      LAYER met4 ;
        RECT 66.330000 197.570000 66.650000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 197.975000 66.650000 198.295000 ;
      LAYER met4 ;
        RECT 66.330000 197.975000 66.650000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 198.380000 66.650000 198.700000 ;
      LAYER met4 ;
        RECT 66.330000 198.380000 66.650000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 198.785000 66.650000 199.105000 ;
      LAYER met4 ;
        RECT 66.330000 198.785000 66.650000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 199.190000 66.650000 199.510000 ;
      LAYER met4 ;
        RECT 66.330000 199.190000 66.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330000 199.595000 66.650000 199.915000 ;
      LAYER met4 ;
        RECT 66.330000 199.595000 66.650000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 175.995000 66.590000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 176.395000 66.590000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 176.795000 66.590000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 177.195000 66.590000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 177.595000 66.590000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 177.995000 66.590000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 178.395000 66.590000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 178.795000 66.590000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 179.195000 66.590000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 179.595000 66.590000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 179.995000 66.590000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 180.395000 66.590000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 180.795000 66.590000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 181.195000 66.590000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 181.595000 66.590000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 181.995000 66.590000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 182.395000 66.590000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 182.795000 66.590000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 183.195000 66.590000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 183.595000 66.590000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 183.995000 66.590000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 184.395000 66.590000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 184.795000 66.590000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 185.195000 66.590000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 185.595000 66.590000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 185.995000 66.590000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 186.395000 66.590000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 186.795000 66.590000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 187.195000 66.590000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 187.595000 66.590000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 187.995000 66.590000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 188.395000 66.590000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 188.795000 66.590000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 189.195000 66.590000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 189.595000 66.590000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 189.995000 66.590000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 190.395000 66.590000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 190.795000 66.590000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 191.195000 66.590000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 191.595000 66.590000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 191.995000 66.590000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 192.395000 66.590000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 192.795000 66.590000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 193.195000 66.590000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 193.595000 66.590000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 193.995000 66.590000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 194.395000 66.590000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.390000 194.795000 66.590000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 25.850000 66.970000 26.170000 ;
      LAYER met4 ;
        RECT 66.650000 25.850000 66.970000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 26.280000 66.970000 26.600000 ;
      LAYER met4 ;
        RECT 66.650000 26.280000 66.970000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 26.710000 66.970000 27.030000 ;
      LAYER met4 ;
        RECT 66.650000 26.710000 66.970000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 27.140000 66.970000 27.460000 ;
      LAYER met4 ;
        RECT 66.650000 27.140000 66.970000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 27.570000 66.970000 27.890000 ;
      LAYER met4 ;
        RECT 66.650000 27.570000 66.970000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 28.000000 66.970000 28.320000 ;
      LAYER met4 ;
        RECT 66.650000 28.000000 66.970000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 28.430000 66.970000 28.750000 ;
      LAYER met4 ;
        RECT 66.650000 28.430000 66.970000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 28.860000 66.970000 29.180000 ;
      LAYER met4 ;
        RECT 66.650000 28.860000 66.970000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 29.290000 66.970000 29.610000 ;
      LAYER met4 ;
        RECT 66.650000 29.290000 66.970000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 29.720000 66.970000 30.040000 ;
      LAYER met4 ;
        RECT 66.650000 29.720000 66.970000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 30.150000 66.970000 30.470000 ;
      LAYER met4 ;
        RECT 66.650000 30.150000 66.970000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 195.140000 67.050000 195.460000 ;
      LAYER met4 ;
        RECT 66.730000 195.140000 67.050000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 195.545000 67.050000 195.865000 ;
      LAYER met4 ;
        RECT 66.730000 195.545000 67.050000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 195.950000 67.050000 196.270000 ;
      LAYER met4 ;
        RECT 66.730000 195.950000 67.050000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 196.355000 67.050000 196.675000 ;
      LAYER met4 ;
        RECT 66.730000 196.355000 67.050000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 196.760000 67.050000 197.080000 ;
      LAYER met4 ;
        RECT 66.730000 196.760000 67.050000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 197.165000 67.050000 197.485000 ;
      LAYER met4 ;
        RECT 66.730000 197.165000 67.050000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 197.570000 67.050000 197.890000 ;
      LAYER met4 ;
        RECT 66.730000 197.570000 67.050000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 197.975000 67.050000 198.295000 ;
      LAYER met4 ;
        RECT 66.730000 197.975000 67.050000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 198.380000 67.050000 198.700000 ;
      LAYER met4 ;
        RECT 66.730000 198.380000 67.050000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 198.785000 67.050000 199.105000 ;
      LAYER met4 ;
        RECT 66.730000 198.785000 67.050000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 199.190000 67.050000 199.510000 ;
      LAYER met4 ;
        RECT 66.730000 199.190000 67.050000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730000 199.595000 67.050000 199.915000 ;
      LAYER met4 ;
        RECT 66.730000 199.595000 67.050000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 175.995000 66.990000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 176.395000 66.990000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 176.795000 66.990000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 177.195000 66.990000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 177.595000 66.990000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 177.995000 66.990000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 178.395000 66.990000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 178.795000 66.990000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 179.195000 66.990000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 179.595000 66.990000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 179.995000 66.990000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 180.395000 66.990000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 180.795000 66.990000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 181.195000 66.990000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 181.595000 66.990000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 181.995000 66.990000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 182.395000 66.990000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 182.795000 66.990000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 183.195000 66.990000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 183.595000 66.990000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 183.995000 66.990000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 184.395000 66.990000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 184.795000 66.990000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 185.195000 66.990000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 185.595000 66.990000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 185.995000 66.990000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 186.395000 66.990000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 186.795000 66.990000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 187.195000 66.990000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 187.595000 66.990000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 187.995000 66.990000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 188.395000 66.990000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 188.795000 66.990000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 189.195000 66.990000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 189.595000 66.990000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 189.995000 66.990000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 190.395000 66.990000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 190.795000 66.990000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 191.195000 66.990000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 191.595000 66.990000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 191.995000 66.990000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 192.395000 66.990000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 192.795000 66.990000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 193.195000 66.990000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 193.595000 66.990000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 193.995000 66.990000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 194.395000 66.990000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.790000 194.795000 66.990000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 25.850000 67.375000 26.170000 ;
      LAYER met4 ;
        RECT 67.055000 25.850000 67.375000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 26.280000 67.375000 26.600000 ;
      LAYER met4 ;
        RECT 67.055000 26.280000 67.375000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 26.710000 67.375000 27.030000 ;
      LAYER met4 ;
        RECT 67.055000 26.710000 67.375000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 27.140000 67.375000 27.460000 ;
      LAYER met4 ;
        RECT 67.055000 27.140000 67.375000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 27.570000 67.375000 27.890000 ;
      LAYER met4 ;
        RECT 67.055000 27.570000 67.375000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 28.000000 67.375000 28.320000 ;
      LAYER met4 ;
        RECT 67.055000 28.000000 67.375000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 28.430000 67.375000 28.750000 ;
      LAYER met4 ;
        RECT 67.055000 28.430000 67.375000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 28.860000 67.375000 29.180000 ;
      LAYER met4 ;
        RECT 67.055000 28.860000 67.375000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 29.290000 67.375000 29.610000 ;
      LAYER met4 ;
        RECT 67.055000 29.290000 67.375000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 29.720000 67.375000 30.040000 ;
      LAYER met4 ;
        RECT 67.055000 29.720000 67.375000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 30.150000 67.375000 30.470000 ;
      LAYER met4 ;
        RECT 67.055000 30.150000 67.375000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 195.140000 67.450000 195.460000 ;
      LAYER met4 ;
        RECT 67.130000 195.140000 67.450000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 195.545000 67.450000 195.865000 ;
      LAYER met4 ;
        RECT 67.130000 195.545000 67.450000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 195.950000 67.450000 196.270000 ;
      LAYER met4 ;
        RECT 67.130000 195.950000 67.450000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 196.355000 67.450000 196.675000 ;
      LAYER met4 ;
        RECT 67.130000 196.355000 67.450000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 196.760000 67.450000 197.080000 ;
      LAYER met4 ;
        RECT 67.130000 196.760000 67.450000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 197.165000 67.450000 197.485000 ;
      LAYER met4 ;
        RECT 67.130000 197.165000 67.450000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 197.570000 67.450000 197.890000 ;
      LAYER met4 ;
        RECT 67.130000 197.570000 67.450000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 197.975000 67.450000 198.295000 ;
      LAYER met4 ;
        RECT 67.130000 197.975000 67.450000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 198.380000 67.450000 198.700000 ;
      LAYER met4 ;
        RECT 67.130000 198.380000 67.450000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 198.785000 67.450000 199.105000 ;
      LAYER met4 ;
        RECT 67.130000 198.785000 67.450000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 199.190000 67.450000 199.510000 ;
      LAYER met4 ;
        RECT 67.130000 199.190000 67.450000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130000 199.595000 67.450000 199.915000 ;
      LAYER met4 ;
        RECT 67.130000 199.595000 67.450000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 175.995000 67.390000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 176.395000 67.390000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 176.795000 67.390000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 177.195000 67.390000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 177.595000 67.390000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 177.995000 67.390000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 178.395000 67.390000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 178.795000 67.390000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 179.195000 67.390000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 179.595000 67.390000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 179.995000 67.390000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 180.395000 67.390000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 180.795000 67.390000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 181.195000 67.390000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 181.595000 67.390000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 181.995000 67.390000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 182.395000 67.390000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 182.795000 67.390000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 183.195000 67.390000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 183.595000 67.390000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 183.995000 67.390000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 184.395000 67.390000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 184.795000 67.390000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 185.195000 67.390000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 185.595000 67.390000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 185.995000 67.390000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 186.395000 67.390000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 186.795000 67.390000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 187.195000 67.390000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 187.595000 67.390000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 187.995000 67.390000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 188.395000 67.390000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 188.795000 67.390000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 189.195000 67.390000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 189.595000 67.390000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 189.995000 67.390000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 190.395000 67.390000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 190.795000 67.390000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 191.195000 67.390000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 191.595000 67.390000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 191.995000 67.390000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 192.395000 67.390000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 192.795000 67.390000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 193.195000 67.390000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 193.595000 67.390000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 193.995000 67.390000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 194.395000 67.390000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.190000 194.795000 67.390000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 25.850000 67.780000 26.170000 ;
      LAYER met4 ;
        RECT 67.460000 25.850000 67.780000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 26.280000 67.780000 26.600000 ;
      LAYER met4 ;
        RECT 67.460000 26.280000 67.780000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 26.710000 67.780000 27.030000 ;
      LAYER met4 ;
        RECT 67.460000 26.710000 67.780000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 27.140000 67.780000 27.460000 ;
      LAYER met4 ;
        RECT 67.460000 27.140000 67.780000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 27.570000 67.780000 27.890000 ;
      LAYER met4 ;
        RECT 67.460000 27.570000 67.780000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 28.000000 67.780000 28.320000 ;
      LAYER met4 ;
        RECT 67.460000 28.000000 67.780000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 28.430000 67.780000 28.750000 ;
      LAYER met4 ;
        RECT 67.460000 28.430000 67.780000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 28.860000 67.780000 29.180000 ;
      LAYER met4 ;
        RECT 67.460000 28.860000 67.780000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 29.290000 67.780000 29.610000 ;
      LAYER met4 ;
        RECT 67.460000 29.290000 67.780000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 29.720000 67.780000 30.040000 ;
      LAYER met4 ;
        RECT 67.460000 29.720000 67.780000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 30.150000 67.780000 30.470000 ;
      LAYER met4 ;
        RECT 67.460000 30.150000 67.780000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 195.140000 67.850000 195.460000 ;
      LAYER met4 ;
        RECT 67.530000 195.140000 67.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 195.545000 67.850000 195.865000 ;
      LAYER met4 ;
        RECT 67.530000 195.545000 67.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 195.950000 67.850000 196.270000 ;
      LAYER met4 ;
        RECT 67.530000 195.950000 67.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 196.355000 67.850000 196.675000 ;
      LAYER met4 ;
        RECT 67.530000 196.355000 67.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 196.760000 67.850000 197.080000 ;
      LAYER met4 ;
        RECT 67.530000 196.760000 67.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 197.165000 67.850000 197.485000 ;
      LAYER met4 ;
        RECT 67.530000 197.165000 67.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 197.570000 67.850000 197.890000 ;
      LAYER met4 ;
        RECT 67.530000 197.570000 67.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 197.975000 67.850000 198.295000 ;
      LAYER met4 ;
        RECT 67.530000 197.975000 67.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 198.380000 67.850000 198.700000 ;
      LAYER met4 ;
        RECT 67.530000 198.380000 67.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 198.785000 67.850000 199.105000 ;
      LAYER met4 ;
        RECT 67.530000 198.785000 67.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 199.190000 67.850000 199.510000 ;
      LAYER met4 ;
        RECT 67.530000 199.190000 67.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530000 199.595000 67.850000 199.915000 ;
      LAYER met4 ;
        RECT 67.530000 199.595000 67.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 175.995000 67.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 176.395000 67.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 176.795000 67.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 177.195000 67.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 177.595000 67.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 177.995000 67.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 178.395000 67.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 178.795000 67.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 179.195000 67.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 179.595000 67.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 179.995000 67.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 180.395000 67.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 180.795000 67.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 181.195000 67.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 181.595000 67.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 181.995000 67.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 182.395000 67.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 182.795000 67.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 183.195000 67.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 183.595000 67.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 183.995000 67.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 184.395000 67.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 184.795000 67.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 185.195000 67.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 185.595000 67.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 185.995000 67.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 186.395000 67.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 186.795000 67.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 187.195000 67.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 187.595000 67.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 187.995000 67.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 188.395000 67.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 188.795000 67.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 189.195000 67.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 189.595000 67.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 189.995000 67.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 190.395000 67.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 190.795000 67.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 191.195000 67.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 191.595000 67.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 191.995000 67.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 192.395000 67.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 192.795000 67.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 193.195000 67.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 193.595000 67.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 193.995000 67.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 194.395000 67.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.590000 194.795000 67.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 25.850000 68.185000 26.170000 ;
      LAYER met4 ;
        RECT 67.865000 25.850000 68.185000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 26.280000 68.185000 26.600000 ;
      LAYER met4 ;
        RECT 67.865000 26.280000 68.185000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 26.710000 68.185000 27.030000 ;
      LAYER met4 ;
        RECT 67.865000 26.710000 68.185000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 27.140000 68.185000 27.460000 ;
      LAYER met4 ;
        RECT 67.865000 27.140000 68.185000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 27.570000 68.185000 27.890000 ;
      LAYER met4 ;
        RECT 67.865000 27.570000 68.185000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 28.000000 68.185000 28.320000 ;
      LAYER met4 ;
        RECT 67.865000 28.000000 68.185000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 28.430000 68.185000 28.750000 ;
      LAYER met4 ;
        RECT 67.865000 28.430000 68.185000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 28.860000 68.185000 29.180000 ;
      LAYER met4 ;
        RECT 67.865000 28.860000 68.185000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 29.290000 68.185000 29.610000 ;
      LAYER met4 ;
        RECT 67.865000 29.290000 68.185000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 29.720000 68.185000 30.040000 ;
      LAYER met4 ;
        RECT 67.865000 29.720000 68.185000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 30.150000 68.185000 30.470000 ;
      LAYER met4 ;
        RECT 67.865000 30.150000 68.185000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 195.140000 68.250000 195.460000 ;
      LAYER met4 ;
        RECT 67.930000 195.140000 68.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 195.545000 68.250000 195.865000 ;
      LAYER met4 ;
        RECT 67.930000 195.545000 68.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 195.950000 68.250000 196.270000 ;
      LAYER met4 ;
        RECT 67.930000 195.950000 68.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 196.355000 68.250000 196.675000 ;
      LAYER met4 ;
        RECT 67.930000 196.355000 68.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 196.760000 68.250000 197.080000 ;
      LAYER met4 ;
        RECT 67.930000 196.760000 68.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 197.165000 68.250000 197.485000 ;
      LAYER met4 ;
        RECT 67.930000 197.165000 68.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 197.570000 68.250000 197.890000 ;
      LAYER met4 ;
        RECT 67.930000 197.570000 68.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 197.975000 68.250000 198.295000 ;
      LAYER met4 ;
        RECT 67.930000 197.975000 68.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 198.380000 68.250000 198.700000 ;
      LAYER met4 ;
        RECT 67.930000 198.380000 68.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 198.785000 68.250000 199.105000 ;
      LAYER met4 ;
        RECT 67.930000 198.785000 68.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 199.190000 68.250000 199.510000 ;
      LAYER met4 ;
        RECT 67.930000 199.190000 68.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930000 199.595000 68.250000 199.915000 ;
      LAYER met4 ;
        RECT 67.930000 199.595000 68.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 175.995000 68.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 176.395000 68.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 176.795000 68.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 177.195000 68.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 177.595000 68.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 177.995000 68.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 178.395000 68.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 178.795000 68.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 179.195000 68.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 179.595000 68.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 179.995000 68.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 180.395000 68.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 180.795000 68.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 181.195000 68.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 181.595000 68.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 181.995000 68.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 182.395000 68.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 182.795000 68.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 183.195000 68.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 183.595000 68.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 183.995000 68.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 184.395000 68.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 184.795000 68.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 185.195000 68.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 185.595000 68.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 185.995000 68.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 186.395000 68.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 186.795000 68.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 187.195000 68.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 187.595000 68.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 187.995000 68.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 188.395000 68.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 188.795000 68.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 189.195000 68.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 189.595000 68.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 189.995000 68.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 190.395000 68.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 190.795000 68.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 191.195000 68.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 191.595000 68.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 191.995000 68.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 192.395000 68.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 192.795000 68.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 193.195000 68.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 193.595000 68.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 193.995000 68.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 194.395000 68.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 194.795000 68.190000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 25.850000 68.590000 26.170000 ;
      LAYER met4 ;
        RECT 68.270000 25.850000 68.590000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 26.280000 68.590000 26.600000 ;
      LAYER met4 ;
        RECT 68.270000 26.280000 68.590000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 26.710000 68.590000 27.030000 ;
      LAYER met4 ;
        RECT 68.270000 26.710000 68.590000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 27.140000 68.590000 27.460000 ;
      LAYER met4 ;
        RECT 68.270000 27.140000 68.590000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 27.570000 68.590000 27.890000 ;
      LAYER met4 ;
        RECT 68.270000 27.570000 68.590000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 28.000000 68.590000 28.320000 ;
      LAYER met4 ;
        RECT 68.270000 28.000000 68.590000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 28.430000 68.590000 28.750000 ;
      LAYER met4 ;
        RECT 68.270000 28.430000 68.590000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 28.860000 68.590000 29.180000 ;
      LAYER met4 ;
        RECT 68.270000 28.860000 68.590000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 29.290000 68.590000 29.610000 ;
      LAYER met4 ;
        RECT 68.270000 29.290000 68.590000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 29.720000 68.590000 30.040000 ;
      LAYER met4 ;
        RECT 68.270000 29.720000 68.590000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 30.150000 68.590000 30.470000 ;
      LAYER met4 ;
        RECT 68.270000 30.150000 68.590000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 195.140000 68.650000 195.460000 ;
      LAYER met4 ;
        RECT 68.330000 195.140000 68.650000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 195.545000 68.650000 195.865000 ;
      LAYER met4 ;
        RECT 68.330000 195.545000 68.650000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 195.950000 68.650000 196.270000 ;
      LAYER met4 ;
        RECT 68.330000 195.950000 68.650000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 196.355000 68.650000 196.675000 ;
      LAYER met4 ;
        RECT 68.330000 196.355000 68.650000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 196.760000 68.650000 197.080000 ;
      LAYER met4 ;
        RECT 68.330000 196.760000 68.650000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 197.165000 68.650000 197.485000 ;
      LAYER met4 ;
        RECT 68.330000 197.165000 68.650000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 197.570000 68.650000 197.890000 ;
      LAYER met4 ;
        RECT 68.330000 197.570000 68.650000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 197.975000 68.650000 198.295000 ;
      LAYER met4 ;
        RECT 68.330000 197.975000 68.650000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 198.380000 68.650000 198.700000 ;
      LAYER met4 ;
        RECT 68.330000 198.380000 68.650000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 198.785000 68.650000 199.105000 ;
      LAYER met4 ;
        RECT 68.330000 198.785000 68.650000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 199.190000 68.650000 199.510000 ;
      LAYER met4 ;
        RECT 68.330000 199.190000 68.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330000 199.595000 68.650000 199.915000 ;
      LAYER met4 ;
        RECT 68.330000 199.595000 68.650000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 175.995000 68.590000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 176.395000 68.590000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 176.795000 68.590000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 177.195000 68.590000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 177.595000 68.590000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 177.995000 68.590000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 178.395000 68.590000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 178.795000 68.590000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 179.195000 68.590000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 179.595000 68.590000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 179.995000 68.590000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 180.395000 68.590000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 180.795000 68.590000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 181.195000 68.590000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 181.595000 68.590000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 181.995000 68.590000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 182.395000 68.590000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 182.795000 68.590000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 183.195000 68.590000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 183.595000 68.590000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 183.995000 68.590000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 184.395000 68.590000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 184.795000 68.590000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 185.195000 68.590000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 185.595000 68.590000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 185.995000 68.590000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 186.395000 68.590000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 186.795000 68.590000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 187.195000 68.590000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 187.595000 68.590000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 187.995000 68.590000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 188.395000 68.590000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 188.795000 68.590000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 189.195000 68.590000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 189.595000 68.590000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 189.995000 68.590000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 190.395000 68.590000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 190.795000 68.590000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 191.195000 68.590000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 191.595000 68.590000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 191.995000 68.590000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 192.395000 68.590000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 192.795000 68.590000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 193.195000 68.590000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 193.595000 68.590000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 193.995000 68.590000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 194.395000 68.590000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.390000 194.795000 68.590000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 25.850000 68.995000 26.170000 ;
      LAYER met4 ;
        RECT 68.675000 25.850000 68.995000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 26.280000 68.995000 26.600000 ;
      LAYER met4 ;
        RECT 68.675000 26.280000 68.995000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 26.710000 68.995000 27.030000 ;
      LAYER met4 ;
        RECT 68.675000 26.710000 68.995000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 27.140000 68.995000 27.460000 ;
      LAYER met4 ;
        RECT 68.675000 27.140000 68.995000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 27.570000 68.995000 27.890000 ;
      LAYER met4 ;
        RECT 68.675000 27.570000 68.995000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 28.000000 68.995000 28.320000 ;
      LAYER met4 ;
        RECT 68.675000 28.000000 68.995000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 28.430000 68.995000 28.750000 ;
      LAYER met4 ;
        RECT 68.675000 28.430000 68.995000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 28.860000 68.995000 29.180000 ;
      LAYER met4 ;
        RECT 68.675000 28.860000 68.995000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 29.290000 68.995000 29.610000 ;
      LAYER met4 ;
        RECT 68.675000 29.290000 68.995000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 29.720000 68.995000 30.040000 ;
      LAYER met4 ;
        RECT 68.675000 29.720000 68.995000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 30.150000 68.995000 30.470000 ;
      LAYER met4 ;
        RECT 68.675000 30.150000 68.995000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 195.140000 69.050000 195.460000 ;
      LAYER met4 ;
        RECT 68.730000 195.140000 69.050000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 195.545000 69.050000 195.865000 ;
      LAYER met4 ;
        RECT 68.730000 195.545000 69.050000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 195.950000 69.050000 196.270000 ;
      LAYER met4 ;
        RECT 68.730000 195.950000 69.050000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 196.355000 69.050000 196.675000 ;
      LAYER met4 ;
        RECT 68.730000 196.355000 69.050000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 196.760000 69.050000 197.080000 ;
      LAYER met4 ;
        RECT 68.730000 196.760000 69.050000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 197.165000 69.050000 197.485000 ;
      LAYER met4 ;
        RECT 68.730000 197.165000 69.050000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 197.570000 69.050000 197.890000 ;
      LAYER met4 ;
        RECT 68.730000 197.570000 69.050000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 197.975000 69.050000 198.295000 ;
      LAYER met4 ;
        RECT 68.730000 197.975000 69.050000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 198.380000 69.050000 198.700000 ;
      LAYER met4 ;
        RECT 68.730000 198.380000 69.050000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 198.785000 69.050000 199.105000 ;
      LAYER met4 ;
        RECT 68.730000 198.785000 69.050000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 199.190000 69.050000 199.510000 ;
      LAYER met4 ;
        RECT 68.730000 199.190000 69.050000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730000 199.595000 69.050000 199.915000 ;
      LAYER met4 ;
        RECT 68.730000 199.595000 69.050000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 175.995000 68.990000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 176.395000 68.990000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 176.795000 68.990000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 177.195000 68.990000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 177.595000 68.990000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 177.995000 68.990000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 178.395000 68.990000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 178.795000 68.990000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 179.195000 68.990000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 179.595000 68.990000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 179.995000 68.990000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 180.395000 68.990000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 180.795000 68.990000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 181.195000 68.990000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 181.595000 68.990000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 181.995000 68.990000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 182.395000 68.990000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 182.795000 68.990000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 183.195000 68.990000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 183.595000 68.990000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 183.995000 68.990000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 184.395000 68.990000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 184.795000 68.990000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 185.195000 68.990000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 185.595000 68.990000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 185.995000 68.990000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 186.395000 68.990000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 186.795000 68.990000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 187.195000 68.990000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 187.595000 68.990000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 187.995000 68.990000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 188.395000 68.990000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 188.795000 68.990000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 189.195000 68.990000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 189.595000 68.990000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 189.995000 68.990000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 190.395000 68.990000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 190.795000 68.990000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 191.195000 68.990000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 191.595000 68.990000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 191.995000 68.990000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 192.395000 68.990000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 192.795000 68.990000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 193.195000 68.990000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 193.595000 68.990000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 193.995000 68.990000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 194.395000 68.990000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.790000 194.795000 68.990000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 25.850000 69.400000 26.170000 ;
      LAYER met4 ;
        RECT 69.080000 25.850000 69.400000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 26.280000 69.400000 26.600000 ;
      LAYER met4 ;
        RECT 69.080000 26.280000 69.400000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 26.710000 69.400000 27.030000 ;
      LAYER met4 ;
        RECT 69.080000 26.710000 69.400000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 27.140000 69.400000 27.460000 ;
      LAYER met4 ;
        RECT 69.080000 27.140000 69.400000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 27.570000 69.400000 27.890000 ;
      LAYER met4 ;
        RECT 69.080000 27.570000 69.400000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 28.000000 69.400000 28.320000 ;
      LAYER met4 ;
        RECT 69.080000 28.000000 69.400000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 28.430000 69.400000 28.750000 ;
      LAYER met4 ;
        RECT 69.080000 28.430000 69.400000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 28.860000 69.400000 29.180000 ;
      LAYER met4 ;
        RECT 69.080000 28.860000 69.400000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 29.290000 69.400000 29.610000 ;
      LAYER met4 ;
        RECT 69.080000 29.290000 69.400000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 29.720000 69.400000 30.040000 ;
      LAYER met4 ;
        RECT 69.080000 29.720000 69.400000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 30.150000 69.400000 30.470000 ;
      LAYER met4 ;
        RECT 69.080000 30.150000 69.400000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 195.140000 69.450000 195.460000 ;
      LAYER met4 ;
        RECT 69.130000 195.140000 69.450000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 195.545000 69.450000 195.865000 ;
      LAYER met4 ;
        RECT 69.130000 195.545000 69.450000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 195.950000 69.450000 196.270000 ;
      LAYER met4 ;
        RECT 69.130000 195.950000 69.450000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 196.355000 69.450000 196.675000 ;
      LAYER met4 ;
        RECT 69.130000 196.355000 69.450000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 196.760000 69.450000 197.080000 ;
      LAYER met4 ;
        RECT 69.130000 196.760000 69.450000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 197.165000 69.450000 197.485000 ;
      LAYER met4 ;
        RECT 69.130000 197.165000 69.450000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 197.570000 69.450000 197.890000 ;
      LAYER met4 ;
        RECT 69.130000 197.570000 69.450000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 197.975000 69.450000 198.295000 ;
      LAYER met4 ;
        RECT 69.130000 197.975000 69.450000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 198.380000 69.450000 198.700000 ;
      LAYER met4 ;
        RECT 69.130000 198.380000 69.450000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 198.785000 69.450000 199.105000 ;
      LAYER met4 ;
        RECT 69.130000 198.785000 69.450000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 199.190000 69.450000 199.510000 ;
      LAYER met4 ;
        RECT 69.130000 199.190000 69.450000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130000 199.595000 69.450000 199.915000 ;
      LAYER met4 ;
        RECT 69.130000 199.595000 69.450000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 175.995000 69.390000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 176.395000 69.390000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 176.795000 69.390000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 177.195000 69.390000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 177.595000 69.390000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 177.995000 69.390000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 178.395000 69.390000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 178.795000 69.390000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 179.195000 69.390000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 179.595000 69.390000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 179.995000 69.390000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 180.395000 69.390000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 180.795000 69.390000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 181.195000 69.390000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 181.595000 69.390000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 181.995000 69.390000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 182.395000 69.390000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 182.795000 69.390000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 183.195000 69.390000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 183.595000 69.390000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 183.995000 69.390000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 184.395000 69.390000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 184.795000 69.390000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 185.195000 69.390000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 185.595000 69.390000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 185.995000 69.390000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 186.395000 69.390000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 186.795000 69.390000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 187.195000 69.390000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 187.595000 69.390000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 187.995000 69.390000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 188.395000 69.390000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 188.795000 69.390000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 189.195000 69.390000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 189.595000 69.390000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 189.995000 69.390000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 190.395000 69.390000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 190.795000 69.390000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 191.195000 69.390000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 191.595000 69.390000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 191.995000 69.390000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 192.395000 69.390000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 192.795000 69.390000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 193.195000 69.390000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 193.595000 69.390000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 193.995000 69.390000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 194.395000 69.390000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 194.795000 69.390000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 25.850000 69.805000 26.170000 ;
      LAYER met4 ;
        RECT 69.485000 25.850000 69.805000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 26.280000 69.805000 26.600000 ;
      LAYER met4 ;
        RECT 69.485000 26.280000 69.805000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 26.710000 69.805000 27.030000 ;
      LAYER met4 ;
        RECT 69.485000 26.710000 69.805000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 27.140000 69.805000 27.460000 ;
      LAYER met4 ;
        RECT 69.485000 27.140000 69.805000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 27.570000 69.805000 27.890000 ;
      LAYER met4 ;
        RECT 69.485000 27.570000 69.805000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 28.000000 69.805000 28.320000 ;
      LAYER met4 ;
        RECT 69.485000 28.000000 69.805000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 28.430000 69.805000 28.750000 ;
      LAYER met4 ;
        RECT 69.485000 28.430000 69.805000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 28.860000 69.805000 29.180000 ;
      LAYER met4 ;
        RECT 69.485000 28.860000 69.805000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 29.290000 69.805000 29.610000 ;
      LAYER met4 ;
        RECT 69.485000 29.290000 69.805000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 29.720000 69.805000 30.040000 ;
      LAYER met4 ;
        RECT 69.485000 29.720000 69.805000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 30.150000 69.805000 30.470000 ;
      LAYER met4 ;
        RECT 69.485000 30.150000 69.805000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 195.140000 69.850000 195.460000 ;
      LAYER met4 ;
        RECT 69.530000 195.140000 69.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 195.545000 69.850000 195.865000 ;
      LAYER met4 ;
        RECT 69.530000 195.545000 69.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 195.950000 69.850000 196.270000 ;
      LAYER met4 ;
        RECT 69.530000 195.950000 69.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 196.355000 69.850000 196.675000 ;
      LAYER met4 ;
        RECT 69.530000 196.355000 69.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 196.760000 69.850000 197.080000 ;
      LAYER met4 ;
        RECT 69.530000 196.760000 69.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 197.165000 69.850000 197.485000 ;
      LAYER met4 ;
        RECT 69.530000 197.165000 69.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 197.570000 69.850000 197.890000 ;
      LAYER met4 ;
        RECT 69.530000 197.570000 69.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 197.975000 69.850000 198.295000 ;
      LAYER met4 ;
        RECT 69.530000 197.975000 69.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 198.380000 69.850000 198.700000 ;
      LAYER met4 ;
        RECT 69.530000 198.380000 69.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 198.785000 69.850000 199.105000 ;
      LAYER met4 ;
        RECT 69.530000 198.785000 69.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 199.190000 69.850000 199.510000 ;
      LAYER met4 ;
        RECT 69.530000 199.190000 69.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530000 199.595000 69.850000 199.915000 ;
      LAYER met4 ;
        RECT 69.530000 199.595000 69.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 175.995000 69.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 176.395000 69.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 176.795000 69.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 177.195000 69.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 177.595000 69.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 177.995000 69.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 178.395000 69.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 178.795000 69.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 179.195000 69.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 179.595000 69.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 179.995000 69.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 180.395000 69.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 180.795000 69.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 181.195000 69.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 181.595000 69.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 181.995000 69.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 182.395000 69.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 182.795000 69.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 183.195000 69.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 183.595000 69.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 183.995000 69.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 184.395000 69.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 184.795000 69.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 185.195000 69.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 185.595000 69.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 185.995000 69.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 186.395000 69.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 186.795000 69.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 187.195000 69.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 187.595000 69.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 187.995000 69.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 188.395000 69.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 188.795000 69.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 189.195000 69.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 189.595000 69.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 189.995000 69.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 190.395000 69.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 190.795000 69.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 191.195000 69.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 191.595000 69.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 191.995000 69.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 192.395000 69.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 192.795000 69.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 193.195000 69.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 193.595000 69.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 193.995000 69.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 194.395000 69.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.590000 194.795000 69.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 25.850000 70.210000 26.170000 ;
      LAYER met4 ;
        RECT 69.890000 25.850000 70.210000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 26.280000 70.210000 26.600000 ;
      LAYER met4 ;
        RECT 69.890000 26.280000 70.210000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 26.710000 70.210000 27.030000 ;
      LAYER met4 ;
        RECT 69.890000 26.710000 70.210000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 27.140000 70.210000 27.460000 ;
      LAYER met4 ;
        RECT 69.890000 27.140000 70.210000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 27.570000 70.210000 27.890000 ;
      LAYER met4 ;
        RECT 69.890000 27.570000 70.210000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 28.000000 70.210000 28.320000 ;
      LAYER met4 ;
        RECT 69.890000 28.000000 70.210000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 28.430000 70.210000 28.750000 ;
      LAYER met4 ;
        RECT 69.890000 28.430000 70.210000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 28.860000 70.210000 29.180000 ;
      LAYER met4 ;
        RECT 69.890000 28.860000 70.210000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 29.290000 70.210000 29.610000 ;
      LAYER met4 ;
        RECT 69.890000 29.290000 70.210000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 29.720000 70.210000 30.040000 ;
      LAYER met4 ;
        RECT 69.890000 29.720000 70.210000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 30.150000 70.210000 30.470000 ;
      LAYER met4 ;
        RECT 69.890000 30.150000 70.210000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 195.140000 70.250000 195.460000 ;
      LAYER met4 ;
        RECT 69.930000 195.140000 70.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 195.545000 70.250000 195.865000 ;
      LAYER met4 ;
        RECT 69.930000 195.545000 70.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 195.950000 70.250000 196.270000 ;
      LAYER met4 ;
        RECT 69.930000 195.950000 70.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 196.355000 70.250000 196.675000 ;
      LAYER met4 ;
        RECT 69.930000 196.355000 70.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 196.760000 70.250000 197.080000 ;
      LAYER met4 ;
        RECT 69.930000 196.760000 70.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 197.165000 70.250000 197.485000 ;
      LAYER met4 ;
        RECT 69.930000 197.165000 70.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 197.570000 70.250000 197.890000 ;
      LAYER met4 ;
        RECT 69.930000 197.570000 70.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 197.975000 70.250000 198.295000 ;
      LAYER met4 ;
        RECT 69.930000 197.975000 70.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 198.380000 70.250000 198.700000 ;
      LAYER met4 ;
        RECT 69.930000 198.380000 70.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 198.785000 70.250000 199.105000 ;
      LAYER met4 ;
        RECT 69.930000 198.785000 70.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 199.190000 70.250000 199.510000 ;
      LAYER met4 ;
        RECT 69.930000 199.190000 70.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930000 199.595000 70.250000 199.915000 ;
      LAYER met4 ;
        RECT 69.930000 199.595000 70.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 175.995000 70.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 176.395000 70.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 176.795000 70.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 177.195000 70.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 177.595000 70.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 177.995000 70.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 178.395000 70.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 178.795000 70.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 179.195000 70.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 179.595000 70.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 179.995000 70.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 180.395000 70.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 180.795000 70.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 181.195000 70.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 181.595000 70.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 181.995000 70.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 182.395000 70.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 182.795000 70.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 183.195000 70.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 183.595000 70.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 183.995000 70.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 184.395000 70.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 184.795000 70.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 185.195000 70.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 185.595000 70.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 185.995000 70.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 186.395000 70.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 186.795000 70.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 187.195000 70.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 187.595000 70.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 187.995000 70.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 188.395000 70.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 188.795000 70.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 189.195000 70.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 189.595000 70.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 189.995000 70.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 190.395000 70.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 190.795000 70.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 191.195000 70.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 191.595000 70.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 191.995000 70.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 192.395000 70.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 192.795000 70.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 193.195000 70.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 193.595000 70.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 193.995000 70.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 194.395000 70.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.990000 194.795000 70.190000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 195.140000 7.345000 195.460000 ;
      LAYER met4 ;
        RECT 7.025000 195.140000 7.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 195.545000 7.345000 195.865000 ;
      LAYER met4 ;
        RECT 7.025000 195.545000 7.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 195.950000 7.345000 196.270000 ;
      LAYER met4 ;
        RECT 7.025000 195.950000 7.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 196.355000 7.345000 196.675000 ;
      LAYER met4 ;
        RECT 7.025000 196.355000 7.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 196.760000 7.345000 197.080000 ;
      LAYER met4 ;
        RECT 7.025000 196.760000 7.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 197.165000 7.345000 197.485000 ;
      LAYER met4 ;
        RECT 7.025000 197.165000 7.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 197.570000 7.345000 197.890000 ;
      LAYER met4 ;
        RECT 7.025000 197.570000 7.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 197.975000 7.345000 198.295000 ;
      LAYER met4 ;
        RECT 7.025000 197.975000 7.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 198.380000 7.345000 198.700000 ;
      LAYER met4 ;
        RECT 7.025000 198.380000 7.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 198.785000 7.345000 199.105000 ;
      LAYER met4 ;
        RECT 7.025000 198.785000 7.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 199.190000 7.345000 199.510000 ;
      LAYER met4 ;
        RECT 7.025000 199.190000 7.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025000 199.595000 7.345000 199.915000 ;
      LAYER met4 ;
        RECT 7.025000 199.595000 7.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 25.850000 7.355000 26.170000 ;
      LAYER met4 ;
        RECT 7.035000 25.850000 7.355000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 26.280000 7.355000 26.600000 ;
      LAYER met4 ;
        RECT 7.035000 26.280000 7.355000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 26.710000 7.355000 27.030000 ;
      LAYER met4 ;
        RECT 7.035000 26.710000 7.355000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 27.140000 7.355000 27.460000 ;
      LAYER met4 ;
        RECT 7.035000 27.140000 7.355000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 27.570000 7.355000 27.890000 ;
      LAYER met4 ;
        RECT 7.035000 27.570000 7.355000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 28.000000 7.355000 28.320000 ;
      LAYER met4 ;
        RECT 7.035000 28.000000 7.355000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 28.430000 7.355000 28.750000 ;
      LAYER met4 ;
        RECT 7.035000 28.430000 7.355000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 28.860000 7.355000 29.180000 ;
      LAYER met4 ;
        RECT 7.035000 28.860000 7.355000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 29.290000 7.355000 29.610000 ;
      LAYER met4 ;
        RECT 7.035000 29.290000 7.355000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 29.720000 7.355000 30.040000 ;
      LAYER met4 ;
        RECT 7.035000 29.720000 7.355000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 30.150000 7.355000 30.470000 ;
      LAYER met4 ;
        RECT 7.035000 30.150000 7.355000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 175.995000 7.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 176.395000 7.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 176.795000 7.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 177.195000 7.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 177.595000 7.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 177.995000 7.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 178.395000 7.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 178.795000 7.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 179.195000 7.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 179.595000 7.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 179.995000 7.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 180.395000 7.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 180.795000 7.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 181.195000 7.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 181.595000 7.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 181.995000 7.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 182.395000 7.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 182.795000 7.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 183.195000 7.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 183.595000 7.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 183.995000 7.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 184.395000 7.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 184.795000 7.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 185.195000 7.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 185.595000 7.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 185.995000 7.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 186.395000 7.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 186.795000 7.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 187.195000 7.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 187.595000 7.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 187.995000 7.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 188.395000 7.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 188.795000 7.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 189.195000 7.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 189.595000 7.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 189.995000 7.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 190.395000 7.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 190.795000 7.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 191.195000 7.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 191.595000 7.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 191.995000 7.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 192.395000 7.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 192.795000 7.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 193.195000 7.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 193.595000 7.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 193.995000 7.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 194.395000 7.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.085000 194.795000 7.285000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 195.140000 7.745000 195.460000 ;
      LAYER met4 ;
        RECT 7.425000 195.140000 7.745000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 195.545000 7.745000 195.865000 ;
      LAYER met4 ;
        RECT 7.425000 195.545000 7.745000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 195.950000 7.745000 196.270000 ;
      LAYER met4 ;
        RECT 7.425000 195.950000 7.745000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 196.355000 7.745000 196.675000 ;
      LAYER met4 ;
        RECT 7.425000 196.355000 7.745000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 196.760000 7.745000 197.080000 ;
      LAYER met4 ;
        RECT 7.425000 196.760000 7.745000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 197.165000 7.745000 197.485000 ;
      LAYER met4 ;
        RECT 7.425000 197.165000 7.745000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 197.570000 7.745000 197.890000 ;
      LAYER met4 ;
        RECT 7.425000 197.570000 7.745000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 197.975000 7.745000 198.295000 ;
      LAYER met4 ;
        RECT 7.425000 197.975000 7.745000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 198.380000 7.745000 198.700000 ;
      LAYER met4 ;
        RECT 7.425000 198.380000 7.745000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 198.785000 7.745000 199.105000 ;
      LAYER met4 ;
        RECT 7.425000 198.785000 7.745000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 199.190000 7.745000 199.510000 ;
      LAYER met4 ;
        RECT 7.425000 199.190000 7.745000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425000 199.595000 7.745000 199.915000 ;
      LAYER met4 ;
        RECT 7.425000 199.595000 7.745000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 25.850000 7.760000 26.170000 ;
      LAYER met4 ;
        RECT 7.440000 25.850000 7.760000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 26.280000 7.760000 26.600000 ;
      LAYER met4 ;
        RECT 7.440000 26.280000 7.760000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 26.710000 7.760000 27.030000 ;
      LAYER met4 ;
        RECT 7.440000 26.710000 7.760000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 27.140000 7.760000 27.460000 ;
      LAYER met4 ;
        RECT 7.440000 27.140000 7.760000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 27.570000 7.760000 27.890000 ;
      LAYER met4 ;
        RECT 7.440000 27.570000 7.760000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 28.000000 7.760000 28.320000 ;
      LAYER met4 ;
        RECT 7.440000 28.000000 7.760000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 28.430000 7.760000 28.750000 ;
      LAYER met4 ;
        RECT 7.440000 28.430000 7.760000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 28.860000 7.760000 29.180000 ;
      LAYER met4 ;
        RECT 7.440000 28.860000 7.760000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 29.290000 7.760000 29.610000 ;
      LAYER met4 ;
        RECT 7.440000 29.290000 7.760000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 29.720000 7.760000 30.040000 ;
      LAYER met4 ;
        RECT 7.440000 29.720000 7.760000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 30.150000 7.760000 30.470000 ;
      LAYER met4 ;
        RECT 7.440000 30.150000 7.760000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 175.995000 7.685000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 176.395000 7.685000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 176.795000 7.685000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 177.195000 7.685000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 177.595000 7.685000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 177.995000 7.685000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 178.395000 7.685000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 178.795000 7.685000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 179.195000 7.685000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 179.595000 7.685000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 179.995000 7.685000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 180.395000 7.685000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 180.795000 7.685000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 181.195000 7.685000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 181.595000 7.685000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 181.995000 7.685000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 182.395000 7.685000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 182.795000 7.685000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 183.195000 7.685000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 183.595000 7.685000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 183.995000 7.685000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 184.395000 7.685000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 184.795000 7.685000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 185.195000 7.685000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 185.595000 7.685000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 185.995000 7.685000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 186.395000 7.685000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 186.795000 7.685000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 187.195000 7.685000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 187.595000 7.685000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 187.995000 7.685000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 188.395000 7.685000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 188.795000 7.685000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 189.195000 7.685000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 189.595000 7.685000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 189.995000 7.685000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 190.395000 7.685000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 190.795000 7.685000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 191.195000 7.685000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 191.595000 7.685000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 191.995000 7.685000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 192.395000 7.685000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 192.795000 7.685000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 193.195000 7.685000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 193.595000 7.685000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 193.995000 7.685000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 194.395000 7.685000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.485000 194.795000 7.685000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 195.140000 8.145000 195.460000 ;
      LAYER met4 ;
        RECT 7.825000 195.140000 8.145000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 195.545000 8.145000 195.865000 ;
      LAYER met4 ;
        RECT 7.825000 195.545000 8.145000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 195.950000 8.145000 196.270000 ;
      LAYER met4 ;
        RECT 7.825000 195.950000 8.145000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 196.355000 8.145000 196.675000 ;
      LAYER met4 ;
        RECT 7.825000 196.355000 8.145000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 196.760000 8.145000 197.080000 ;
      LAYER met4 ;
        RECT 7.825000 196.760000 8.145000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 197.165000 8.145000 197.485000 ;
      LAYER met4 ;
        RECT 7.825000 197.165000 8.145000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 197.570000 8.145000 197.890000 ;
      LAYER met4 ;
        RECT 7.825000 197.570000 8.145000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 197.975000 8.145000 198.295000 ;
      LAYER met4 ;
        RECT 7.825000 197.975000 8.145000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 198.380000 8.145000 198.700000 ;
      LAYER met4 ;
        RECT 7.825000 198.380000 8.145000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 198.785000 8.145000 199.105000 ;
      LAYER met4 ;
        RECT 7.825000 198.785000 8.145000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 199.190000 8.145000 199.510000 ;
      LAYER met4 ;
        RECT 7.825000 199.190000 8.145000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825000 199.595000 8.145000 199.915000 ;
      LAYER met4 ;
        RECT 7.825000 199.595000 8.145000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 25.850000 8.165000 26.170000 ;
      LAYER met4 ;
        RECT 7.845000 25.850000 8.165000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 26.280000 8.165000 26.600000 ;
      LAYER met4 ;
        RECT 7.845000 26.280000 8.165000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 26.710000 8.165000 27.030000 ;
      LAYER met4 ;
        RECT 7.845000 26.710000 8.165000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 27.140000 8.165000 27.460000 ;
      LAYER met4 ;
        RECT 7.845000 27.140000 8.165000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 27.570000 8.165000 27.890000 ;
      LAYER met4 ;
        RECT 7.845000 27.570000 8.165000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 28.000000 8.165000 28.320000 ;
      LAYER met4 ;
        RECT 7.845000 28.000000 8.165000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 28.430000 8.165000 28.750000 ;
      LAYER met4 ;
        RECT 7.845000 28.430000 8.165000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 28.860000 8.165000 29.180000 ;
      LAYER met4 ;
        RECT 7.845000 28.860000 8.165000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 29.290000 8.165000 29.610000 ;
      LAYER met4 ;
        RECT 7.845000 29.290000 8.165000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 29.720000 8.165000 30.040000 ;
      LAYER met4 ;
        RECT 7.845000 29.720000 8.165000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 30.150000 8.165000 30.470000 ;
      LAYER met4 ;
        RECT 7.845000 30.150000 8.165000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 175.995000 8.085000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 176.395000 8.085000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 176.795000 8.085000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 177.195000 8.085000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 177.595000 8.085000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 177.995000 8.085000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 178.395000 8.085000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 178.795000 8.085000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 179.195000 8.085000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 179.595000 8.085000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 179.995000 8.085000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 180.395000 8.085000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 180.795000 8.085000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 181.195000 8.085000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 181.595000 8.085000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 181.995000 8.085000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 182.395000 8.085000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 182.795000 8.085000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 183.195000 8.085000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 183.595000 8.085000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 183.995000 8.085000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 184.395000 8.085000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 184.795000 8.085000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 185.195000 8.085000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 185.595000 8.085000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 185.995000 8.085000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 186.395000 8.085000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 186.795000 8.085000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 187.195000 8.085000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 187.595000 8.085000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 187.995000 8.085000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 188.395000 8.085000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 188.795000 8.085000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 189.195000 8.085000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 189.595000 8.085000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 189.995000 8.085000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 190.395000 8.085000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 190.795000 8.085000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 191.195000 8.085000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 191.595000 8.085000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 191.995000 8.085000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 192.395000 8.085000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 192.795000 8.085000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 193.195000 8.085000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 193.595000 8.085000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 193.995000 8.085000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 194.395000 8.085000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 194.795000 8.085000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 25.850000 70.615000 26.170000 ;
      LAYER met4 ;
        RECT 70.295000 25.850000 70.615000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 26.280000 70.615000 26.600000 ;
      LAYER met4 ;
        RECT 70.295000 26.280000 70.615000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 26.710000 70.615000 27.030000 ;
      LAYER met4 ;
        RECT 70.295000 26.710000 70.615000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 27.140000 70.615000 27.460000 ;
      LAYER met4 ;
        RECT 70.295000 27.140000 70.615000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 27.570000 70.615000 27.890000 ;
      LAYER met4 ;
        RECT 70.295000 27.570000 70.615000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 28.000000 70.615000 28.320000 ;
      LAYER met4 ;
        RECT 70.295000 28.000000 70.615000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 28.430000 70.615000 28.750000 ;
      LAYER met4 ;
        RECT 70.295000 28.430000 70.615000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 28.860000 70.615000 29.180000 ;
      LAYER met4 ;
        RECT 70.295000 28.860000 70.615000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 29.290000 70.615000 29.610000 ;
      LAYER met4 ;
        RECT 70.295000 29.290000 70.615000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 29.720000 70.615000 30.040000 ;
      LAYER met4 ;
        RECT 70.295000 29.720000 70.615000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 30.150000 70.615000 30.470000 ;
      LAYER met4 ;
        RECT 70.295000 30.150000 70.615000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 195.140000 70.650000 195.460000 ;
      LAYER met4 ;
        RECT 70.330000 195.140000 70.650000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 195.545000 70.650000 195.865000 ;
      LAYER met4 ;
        RECT 70.330000 195.545000 70.650000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 195.950000 70.650000 196.270000 ;
      LAYER met4 ;
        RECT 70.330000 195.950000 70.650000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 196.355000 70.650000 196.675000 ;
      LAYER met4 ;
        RECT 70.330000 196.355000 70.650000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 196.760000 70.650000 197.080000 ;
      LAYER met4 ;
        RECT 70.330000 196.760000 70.650000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 197.165000 70.650000 197.485000 ;
      LAYER met4 ;
        RECT 70.330000 197.165000 70.650000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 197.570000 70.650000 197.890000 ;
      LAYER met4 ;
        RECT 70.330000 197.570000 70.650000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 197.975000 70.650000 198.295000 ;
      LAYER met4 ;
        RECT 70.330000 197.975000 70.650000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 198.380000 70.650000 198.700000 ;
      LAYER met4 ;
        RECT 70.330000 198.380000 70.650000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 198.785000 70.650000 199.105000 ;
      LAYER met4 ;
        RECT 70.330000 198.785000 70.650000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 199.190000 70.650000 199.510000 ;
      LAYER met4 ;
        RECT 70.330000 199.190000 70.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330000 199.595000 70.650000 199.915000 ;
      LAYER met4 ;
        RECT 70.330000 199.595000 70.650000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 175.995000 70.590000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 176.395000 70.590000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 176.795000 70.590000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 177.195000 70.590000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 177.595000 70.590000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 177.995000 70.590000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 178.395000 70.590000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 178.795000 70.590000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 179.195000 70.590000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 179.595000 70.590000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 179.995000 70.590000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 180.395000 70.590000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 180.795000 70.590000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 181.195000 70.590000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 181.595000 70.590000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 181.995000 70.590000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 182.395000 70.590000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 182.795000 70.590000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 183.195000 70.590000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 183.595000 70.590000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 183.995000 70.590000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 184.395000 70.590000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 184.795000 70.590000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 185.195000 70.590000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 185.595000 70.590000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 185.995000 70.590000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 186.395000 70.590000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 186.795000 70.590000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 187.195000 70.590000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 187.595000 70.590000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 187.995000 70.590000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 188.395000 70.590000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 188.795000 70.590000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 189.195000 70.590000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 189.595000 70.590000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 189.995000 70.590000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 190.395000 70.590000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 190.795000 70.590000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 191.195000 70.590000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 191.595000 70.590000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 191.995000 70.590000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 192.395000 70.590000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 192.795000 70.590000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 193.195000 70.590000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 193.595000 70.590000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 193.995000 70.590000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 194.395000 70.590000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 194.795000 70.590000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 25.850000 71.020000 26.170000 ;
      LAYER met4 ;
        RECT 70.700000 25.850000 71.020000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 26.280000 71.020000 26.600000 ;
      LAYER met4 ;
        RECT 70.700000 26.280000 71.020000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 26.710000 71.020000 27.030000 ;
      LAYER met4 ;
        RECT 70.700000 26.710000 71.020000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 27.140000 71.020000 27.460000 ;
      LAYER met4 ;
        RECT 70.700000 27.140000 71.020000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 27.570000 71.020000 27.890000 ;
      LAYER met4 ;
        RECT 70.700000 27.570000 71.020000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 28.000000 71.020000 28.320000 ;
      LAYER met4 ;
        RECT 70.700000 28.000000 71.020000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 28.430000 71.020000 28.750000 ;
      LAYER met4 ;
        RECT 70.700000 28.430000 71.020000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 28.860000 71.020000 29.180000 ;
      LAYER met4 ;
        RECT 70.700000 28.860000 71.020000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 29.290000 71.020000 29.610000 ;
      LAYER met4 ;
        RECT 70.700000 29.290000 71.020000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 29.720000 71.020000 30.040000 ;
      LAYER met4 ;
        RECT 70.700000 29.720000 71.020000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 30.150000 71.020000 30.470000 ;
      LAYER met4 ;
        RECT 70.700000 30.150000 71.020000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 195.140000 71.050000 195.460000 ;
      LAYER met4 ;
        RECT 70.730000 195.140000 71.050000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 195.545000 71.050000 195.865000 ;
      LAYER met4 ;
        RECT 70.730000 195.545000 71.050000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 195.950000 71.050000 196.270000 ;
      LAYER met4 ;
        RECT 70.730000 195.950000 71.050000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 196.355000 71.050000 196.675000 ;
      LAYER met4 ;
        RECT 70.730000 196.355000 71.050000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 196.760000 71.050000 197.080000 ;
      LAYER met4 ;
        RECT 70.730000 196.760000 71.050000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 197.165000 71.050000 197.485000 ;
      LAYER met4 ;
        RECT 70.730000 197.165000 71.050000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 197.570000 71.050000 197.890000 ;
      LAYER met4 ;
        RECT 70.730000 197.570000 71.050000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 197.975000 71.050000 198.295000 ;
      LAYER met4 ;
        RECT 70.730000 197.975000 71.050000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 198.380000 71.050000 198.700000 ;
      LAYER met4 ;
        RECT 70.730000 198.380000 71.050000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 198.785000 71.050000 199.105000 ;
      LAYER met4 ;
        RECT 70.730000 198.785000 71.050000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 199.190000 71.050000 199.510000 ;
      LAYER met4 ;
        RECT 70.730000 199.190000 71.050000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730000 199.595000 71.050000 199.915000 ;
      LAYER met4 ;
        RECT 70.730000 199.595000 71.050000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 175.995000 70.990000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 176.395000 70.990000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 176.795000 70.990000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 177.195000 70.990000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 177.595000 70.990000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 177.995000 70.990000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 178.395000 70.990000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 178.795000 70.990000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 179.195000 70.990000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 179.595000 70.990000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 179.995000 70.990000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 180.395000 70.990000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 180.795000 70.990000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 181.195000 70.990000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 181.595000 70.990000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 181.995000 70.990000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 182.395000 70.990000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 182.795000 70.990000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 183.195000 70.990000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 183.595000 70.990000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 183.995000 70.990000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 184.395000 70.990000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 184.795000 70.990000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 185.195000 70.990000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 185.595000 70.990000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 185.995000 70.990000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 186.395000 70.990000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 186.795000 70.990000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 187.195000 70.990000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 187.595000 70.990000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 187.995000 70.990000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 188.395000 70.990000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 188.795000 70.990000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 189.195000 70.990000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 189.595000 70.990000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 189.995000 70.990000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 190.395000 70.990000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 190.795000 70.990000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 191.195000 70.990000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 191.595000 70.990000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 191.995000 70.990000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 192.395000 70.990000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 192.795000 70.990000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 193.195000 70.990000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 193.595000 70.990000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 193.995000 70.990000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 194.395000 70.990000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.790000 194.795000 70.990000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 25.850000 71.425000 26.170000 ;
      LAYER met4 ;
        RECT 71.105000 25.850000 71.425000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 26.280000 71.425000 26.600000 ;
      LAYER met4 ;
        RECT 71.105000 26.280000 71.425000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 26.710000 71.425000 27.030000 ;
      LAYER met4 ;
        RECT 71.105000 26.710000 71.425000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 27.140000 71.425000 27.460000 ;
      LAYER met4 ;
        RECT 71.105000 27.140000 71.425000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 27.570000 71.425000 27.890000 ;
      LAYER met4 ;
        RECT 71.105000 27.570000 71.425000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 28.000000 71.425000 28.320000 ;
      LAYER met4 ;
        RECT 71.105000 28.000000 71.425000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 28.430000 71.425000 28.750000 ;
      LAYER met4 ;
        RECT 71.105000 28.430000 71.425000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 28.860000 71.425000 29.180000 ;
      LAYER met4 ;
        RECT 71.105000 28.860000 71.425000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 29.290000 71.425000 29.610000 ;
      LAYER met4 ;
        RECT 71.105000 29.290000 71.425000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 29.720000 71.425000 30.040000 ;
      LAYER met4 ;
        RECT 71.105000 29.720000 71.425000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 30.150000 71.425000 30.470000 ;
      LAYER met4 ;
        RECT 71.105000 30.150000 71.425000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 195.140000 71.450000 195.460000 ;
      LAYER met4 ;
        RECT 71.130000 195.140000 71.450000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 195.545000 71.450000 195.865000 ;
      LAYER met4 ;
        RECT 71.130000 195.545000 71.450000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 195.950000 71.450000 196.270000 ;
      LAYER met4 ;
        RECT 71.130000 195.950000 71.450000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 196.355000 71.450000 196.675000 ;
      LAYER met4 ;
        RECT 71.130000 196.355000 71.450000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 196.760000 71.450000 197.080000 ;
      LAYER met4 ;
        RECT 71.130000 196.760000 71.450000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 197.165000 71.450000 197.485000 ;
      LAYER met4 ;
        RECT 71.130000 197.165000 71.450000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 197.570000 71.450000 197.890000 ;
      LAYER met4 ;
        RECT 71.130000 197.570000 71.450000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 197.975000 71.450000 198.295000 ;
      LAYER met4 ;
        RECT 71.130000 197.975000 71.450000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 198.380000 71.450000 198.700000 ;
      LAYER met4 ;
        RECT 71.130000 198.380000 71.450000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 198.785000 71.450000 199.105000 ;
      LAYER met4 ;
        RECT 71.130000 198.785000 71.450000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 199.190000 71.450000 199.510000 ;
      LAYER met4 ;
        RECT 71.130000 199.190000 71.450000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130000 199.595000 71.450000 199.915000 ;
      LAYER met4 ;
        RECT 71.130000 199.595000 71.450000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 175.995000 71.390000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 176.395000 71.390000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 176.795000 71.390000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 177.195000 71.390000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 177.595000 71.390000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 177.995000 71.390000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 178.395000 71.390000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 178.795000 71.390000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 179.195000 71.390000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 179.595000 71.390000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 179.995000 71.390000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 180.395000 71.390000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 180.795000 71.390000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 181.195000 71.390000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 181.595000 71.390000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 181.995000 71.390000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 182.395000 71.390000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 182.795000 71.390000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 183.195000 71.390000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 183.595000 71.390000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 183.995000 71.390000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 184.395000 71.390000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 184.795000 71.390000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 185.195000 71.390000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 185.595000 71.390000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 185.995000 71.390000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 186.395000 71.390000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 186.795000 71.390000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 187.195000 71.390000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 187.595000 71.390000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 187.995000 71.390000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 188.395000 71.390000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 188.795000 71.390000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 189.195000 71.390000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 189.595000 71.390000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 189.995000 71.390000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 190.395000 71.390000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 190.795000 71.390000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 191.195000 71.390000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 191.595000 71.390000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 191.995000 71.390000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 192.395000 71.390000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 192.795000 71.390000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 193.195000 71.390000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 193.595000 71.390000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 193.995000 71.390000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 194.395000 71.390000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.190000 194.795000 71.390000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 25.850000 71.830000 26.170000 ;
      LAYER met4 ;
        RECT 71.510000 25.850000 71.830000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 26.280000 71.830000 26.600000 ;
      LAYER met4 ;
        RECT 71.510000 26.280000 71.830000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 26.710000 71.830000 27.030000 ;
      LAYER met4 ;
        RECT 71.510000 26.710000 71.830000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 27.140000 71.830000 27.460000 ;
      LAYER met4 ;
        RECT 71.510000 27.140000 71.830000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 27.570000 71.830000 27.890000 ;
      LAYER met4 ;
        RECT 71.510000 27.570000 71.830000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 28.000000 71.830000 28.320000 ;
      LAYER met4 ;
        RECT 71.510000 28.000000 71.830000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 28.430000 71.830000 28.750000 ;
      LAYER met4 ;
        RECT 71.510000 28.430000 71.830000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 28.860000 71.830000 29.180000 ;
      LAYER met4 ;
        RECT 71.510000 28.860000 71.830000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 29.290000 71.830000 29.610000 ;
      LAYER met4 ;
        RECT 71.510000 29.290000 71.830000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 29.720000 71.830000 30.040000 ;
      LAYER met4 ;
        RECT 71.510000 29.720000 71.830000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 30.150000 71.830000 30.470000 ;
      LAYER met4 ;
        RECT 71.510000 30.150000 71.830000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 195.140000 71.850000 195.460000 ;
      LAYER met4 ;
        RECT 71.530000 195.140000 71.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 195.545000 71.850000 195.865000 ;
      LAYER met4 ;
        RECT 71.530000 195.545000 71.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 195.950000 71.850000 196.270000 ;
      LAYER met4 ;
        RECT 71.530000 195.950000 71.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 196.355000 71.850000 196.675000 ;
      LAYER met4 ;
        RECT 71.530000 196.355000 71.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 196.760000 71.850000 197.080000 ;
      LAYER met4 ;
        RECT 71.530000 196.760000 71.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 197.165000 71.850000 197.485000 ;
      LAYER met4 ;
        RECT 71.530000 197.165000 71.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 197.570000 71.850000 197.890000 ;
      LAYER met4 ;
        RECT 71.530000 197.570000 71.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 197.975000 71.850000 198.295000 ;
      LAYER met4 ;
        RECT 71.530000 197.975000 71.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 198.380000 71.850000 198.700000 ;
      LAYER met4 ;
        RECT 71.530000 198.380000 71.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 198.785000 71.850000 199.105000 ;
      LAYER met4 ;
        RECT 71.530000 198.785000 71.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 199.190000 71.850000 199.510000 ;
      LAYER met4 ;
        RECT 71.530000 199.190000 71.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530000 199.595000 71.850000 199.915000 ;
      LAYER met4 ;
        RECT 71.530000 199.595000 71.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 175.995000 71.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 176.395000 71.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 176.795000 71.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 177.195000 71.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 177.595000 71.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 177.995000 71.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 178.395000 71.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 178.795000 71.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 179.195000 71.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 179.595000 71.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 179.995000 71.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 180.395000 71.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 180.795000 71.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 181.195000 71.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 181.595000 71.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 181.995000 71.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 182.395000 71.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 182.795000 71.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 183.195000 71.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 183.595000 71.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 183.995000 71.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 184.395000 71.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 184.795000 71.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 185.195000 71.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 185.595000 71.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 185.995000 71.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 186.395000 71.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 186.795000 71.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 187.195000 71.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 187.595000 71.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 187.995000 71.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 188.395000 71.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 188.795000 71.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 189.195000 71.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 189.595000 71.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 189.995000 71.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 190.395000 71.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 190.795000 71.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 191.195000 71.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 191.595000 71.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 191.995000 71.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 192.395000 71.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 192.795000 71.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 193.195000 71.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 193.595000 71.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 193.995000 71.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 194.395000 71.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 194.795000 71.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 25.850000 72.235000 26.170000 ;
      LAYER met4 ;
        RECT 71.915000 25.850000 72.235000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 26.280000 72.235000 26.600000 ;
      LAYER met4 ;
        RECT 71.915000 26.280000 72.235000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 26.710000 72.235000 27.030000 ;
      LAYER met4 ;
        RECT 71.915000 26.710000 72.235000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 27.140000 72.235000 27.460000 ;
      LAYER met4 ;
        RECT 71.915000 27.140000 72.235000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 27.570000 72.235000 27.890000 ;
      LAYER met4 ;
        RECT 71.915000 27.570000 72.235000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 28.000000 72.235000 28.320000 ;
      LAYER met4 ;
        RECT 71.915000 28.000000 72.235000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 28.430000 72.235000 28.750000 ;
      LAYER met4 ;
        RECT 71.915000 28.430000 72.235000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 28.860000 72.235000 29.180000 ;
      LAYER met4 ;
        RECT 71.915000 28.860000 72.235000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 29.290000 72.235000 29.610000 ;
      LAYER met4 ;
        RECT 71.915000 29.290000 72.235000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 29.720000 72.235000 30.040000 ;
      LAYER met4 ;
        RECT 71.915000 29.720000 72.235000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 30.150000 72.235000 30.470000 ;
      LAYER met4 ;
        RECT 71.915000 30.150000 72.235000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 195.140000 72.250000 195.460000 ;
      LAYER met4 ;
        RECT 71.930000 195.140000 72.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 195.545000 72.250000 195.865000 ;
      LAYER met4 ;
        RECT 71.930000 195.545000 72.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 195.950000 72.250000 196.270000 ;
      LAYER met4 ;
        RECT 71.930000 195.950000 72.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 196.355000 72.250000 196.675000 ;
      LAYER met4 ;
        RECT 71.930000 196.355000 72.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 196.760000 72.250000 197.080000 ;
      LAYER met4 ;
        RECT 71.930000 196.760000 72.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 197.165000 72.250000 197.485000 ;
      LAYER met4 ;
        RECT 71.930000 197.165000 72.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 197.570000 72.250000 197.890000 ;
      LAYER met4 ;
        RECT 71.930000 197.570000 72.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 197.975000 72.250000 198.295000 ;
      LAYER met4 ;
        RECT 71.930000 197.975000 72.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 198.380000 72.250000 198.700000 ;
      LAYER met4 ;
        RECT 71.930000 198.380000 72.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 198.785000 72.250000 199.105000 ;
      LAYER met4 ;
        RECT 71.930000 198.785000 72.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 199.190000 72.250000 199.510000 ;
      LAYER met4 ;
        RECT 71.930000 199.190000 72.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930000 199.595000 72.250000 199.915000 ;
      LAYER met4 ;
        RECT 71.930000 199.595000 72.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 175.995000 72.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 176.395000 72.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 176.795000 72.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 177.195000 72.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 177.595000 72.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 177.995000 72.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 178.395000 72.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 178.795000 72.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 179.195000 72.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 179.595000 72.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 179.995000 72.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 180.395000 72.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 180.795000 72.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 181.195000 72.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 181.595000 72.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 181.995000 72.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 182.395000 72.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 182.795000 72.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 183.195000 72.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 183.595000 72.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 183.995000 72.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 184.395000 72.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 184.795000 72.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 185.195000 72.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 185.595000 72.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 185.995000 72.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 186.395000 72.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 186.795000 72.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 187.195000 72.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 187.595000 72.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 187.995000 72.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 188.395000 72.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 188.795000 72.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 189.195000 72.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 189.595000 72.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 189.995000 72.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 190.395000 72.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 190.795000 72.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 191.195000 72.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 191.595000 72.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 191.995000 72.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 192.395000 72.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 192.795000 72.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 193.195000 72.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 193.595000 72.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 193.995000 72.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 194.395000 72.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.990000 194.795000 72.190000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 25.850000 72.640000 26.170000 ;
      LAYER met4 ;
        RECT 72.320000 25.850000 72.640000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 26.280000 72.640000 26.600000 ;
      LAYER met4 ;
        RECT 72.320000 26.280000 72.640000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 26.710000 72.640000 27.030000 ;
      LAYER met4 ;
        RECT 72.320000 26.710000 72.640000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 27.140000 72.640000 27.460000 ;
      LAYER met4 ;
        RECT 72.320000 27.140000 72.640000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 27.570000 72.640000 27.890000 ;
      LAYER met4 ;
        RECT 72.320000 27.570000 72.640000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 28.000000 72.640000 28.320000 ;
      LAYER met4 ;
        RECT 72.320000 28.000000 72.640000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 28.430000 72.640000 28.750000 ;
      LAYER met4 ;
        RECT 72.320000 28.430000 72.640000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 28.860000 72.640000 29.180000 ;
      LAYER met4 ;
        RECT 72.320000 28.860000 72.640000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 29.290000 72.640000 29.610000 ;
      LAYER met4 ;
        RECT 72.320000 29.290000 72.640000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 29.720000 72.640000 30.040000 ;
      LAYER met4 ;
        RECT 72.320000 29.720000 72.640000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 30.150000 72.640000 30.470000 ;
      LAYER met4 ;
        RECT 72.320000 30.150000 72.640000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 195.140000 72.650000 195.460000 ;
      LAYER met4 ;
        RECT 72.330000 195.140000 72.650000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 195.545000 72.650000 195.865000 ;
      LAYER met4 ;
        RECT 72.330000 195.545000 72.650000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 195.950000 72.650000 196.270000 ;
      LAYER met4 ;
        RECT 72.330000 195.950000 72.650000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 196.355000 72.650000 196.675000 ;
      LAYER met4 ;
        RECT 72.330000 196.355000 72.650000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 196.760000 72.650000 197.080000 ;
      LAYER met4 ;
        RECT 72.330000 196.760000 72.650000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 197.165000 72.650000 197.485000 ;
      LAYER met4 ;
        RECT 72.330000 197.165000 72.650000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 197.570000 72.650000 197.890000 ;
      LAYER met4 ;
        RECT 72.330000 197.570000 72.650000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 197.975000 72.650000 198.295000 ;
      LAYER met4 ;
        RECT 72.330000 197.975000 72.650000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 198.380000 72.650000 198.700000 ;
      LAYER met4 ;
        RECT 72.330000 198.380000 72.650000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 198.785000 72.650000 199.105000 ;
      LAYER met4 ;
        RECT 72.330000 198.785000 72.650000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 199.190000 72.650000 199.510000 ;
      LAYER met4 ;
        RECT 72.330000 199.190000 72.650000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 199.595000 72.650000 199.915000 ;
      LAYER met4 ;
        RECT 72.330000 199.595000 72.650000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 175.995000 72.590000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 176.395000 72.590000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 176.795000 72.590000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 177.195000 72.590000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 177.595000 72.590000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 177.995000 72.590000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 178.395000 72.590000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 178.795000 72.590000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 179.195000 72.590000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 179.595000 72.590000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 179.995000 72.590000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 180.395000 72.590000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 180.795000 72.590000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 181.195000 72.590000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 181.595000 72.590000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 181.995000 72.590000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 182.395000 72.590000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 182.795000 72.590000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 183.195000 72.590000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 183.595000 72.590000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 183.995000 72.590000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 184.395000 72.590000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 184.795000 72.590000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 185.195000 72.590000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 185.595000 72.590000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 185.995000 72.590000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 186.395000 72.590000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 186.795000 72.590000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 187.195000 72.590000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 187.595000 72.590000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 187.995000 72.590000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 188.395000 72.590000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 188.795000 72.590000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 189.195000 72.590000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 189.595000 72.590000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 189.995000 72.590000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 190.395000 72.590000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 190.795000 72.590000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 191.195000 72.590000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 191.595000 72.590000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 191.995000 72.590000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 192.395000 72.590000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 192.795000 72.590000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 193.195000 72.590000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 193.595000 72.590000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 193.995000 72.590000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 194.395000 72.590000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390000 194.795000 72.590000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 25.850000 73.045000 26.170000 ;
      LAYER met4 ;
        RECT 72.725000 25.850000 73.045000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 26.280000 73.045000 26.600000 ;
      LAYER met4 ;
        RECT 72.725000 26.280000 73.045000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 26.710000 73.045000 27.030000 ;
      LAYER met4 ;
        RECT 72.725000 26.710000 73.045000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 27.140000 73.045000 27.460000 ;
      LAYER met4 ;
        RECT 72.725000 27.140000 73.045000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 27.570000 73.045000 27.890000 ;
      LAYER met4 ;
        RECT 72.725000 27.570000 73.045000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 28.000000 73.045000 28.320000 ;
      LAYER met4 ;
        RECT 72.725000 28.000000 73.045000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 28.430000 73.045000 28.750000 ;
      LAYER met4 ;
        RECT 72.725000 28.430000 73.045000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 28.860000 73.045000 29.180000 ;
      LAYER met4 ;
        RECT 72.725000 28.860000 73.045000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 29.290000 73.045000 29.610000 ;
      LAYER met4 ;
        RECT 72.725000 29.290000 73.045000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 29.720000 73.045000 30.040000 ;
      LAYER met4 ;
        RECT 72.725000 29.720000 73.045000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 30.150000 73.045000 30.470000 ;
      LAYER met4 ;
        RECT 72.725000 30.150000 73.045000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 195.140000 73.050000 195.460000 ;
      LAYER met4 ;
        RECT 72.730000 195.140000 73.050000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 195.545000 73.050000 195.865000 ;
      LAYER met4 ;
        RECT 72.730000 195.545000 73.050000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 195.950000 73.050000 196.270000 ;
      LAYER met4 ;
        RECT 72.730000 195.950000 73.050000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 196.355000 73.050000 196.675000 ;
      LAYER met4 ;
        RECT 72.730000 196.355000 73.050000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 196.760000 73.050000 197.080000 ;
      LAYER met4 ;
        RECT 72.730000 196.760000 73.050000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 197.165000 73.050000 197.485000 ;
      LAYER met4 ;
        RECT 72.730000 197.165000 73.050000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 197.570000 73.050000 197.890000 ;
      LAYER met4 ;
        RECT 72.730000 197.570000 73.050000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 197.975000 73.050000 198.295000 ;
      LAYER met4 ;
        RECT 72.730000 197.975000 73.050000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 198.380000 73.050000 198.700000 ;
      LAYER met4 ;
        RECT 72.730000 198.380000 73.050000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 198.785000 73.050000 199.105000 ;
      LAYER met4 ;
        RECT 72.730000 198.785000 73.050000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 199.190000 73.050000 199.510000 ;
      LAYER met4 ;
        RECT 72.730000 199.190000 73.050000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 199.595000 73.050000 199.915000 ;
      LAYER met4 ;
        RECT 72.730000 199.595000 73.050000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 175.995000 72.990000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 176.395000 72.990000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 176.795000 72.990000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 177.195000 72.990000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 177.595000 72.990000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 177.995000 72.990000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 178.395000 72.990000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 178.795000 72.990000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 179.195000 72.990000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 179.595000 72.990000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 179.995000 72.990000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 180.395000 72.990000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 180.795000 72.990000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 181.195000 72.990000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 181.595000 72.990000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 181.995000 72.990000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 182.395000 72.990000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 182.795000 72.990000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 183.195000 72.990000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 183.595000 72.990000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 183.995000 72.990000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 184.395000 72.990000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 184.795000 72.990000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 185.195000 72.990000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 185.595000 72.990000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 185.995000 72.990000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 186.395000 72.990000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 186.795000 72.990000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 187.195000 72.990000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 187.595000 72.990000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 187.995000 72.990000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 188.395000 72.990000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 188.795000 72.990000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 189.195000 72.990000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 189.595000 72.990000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 189.995000 72.990000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 190.395000 72.990000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 190.795000 72.990000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 191.195000 72.990000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 191.595000 72.990000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 191.995000 72.990000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 192.395000 72.990000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 192.795000 72.990000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 193.195000 72.990000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 193.595000 72.990000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 193.995000 72.990000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 194.395000 72.990000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790000 194.795000 72.990000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 195.140000 73.450000 195.460000 ;
      LAYER met4 ;
        RECT 73.130000 195.140000 73.450000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 195.545000 73.450000 195.865000 ;
      LAYER met4 ;
        RECT 73.130000 195.545000 73.450000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 195.950000 73.450000 196.270000 ;
      LAYER met4 ;
        RECT 73.130000 195.950000 73.450000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 196.355000 73.450000 196.675000 ;
      LAYER met4 ;
        RECT 73.130000 196.355000 73.450000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 196.760000 73.450000 197.080000 ;
      LAYER met4 ;
        RECT 73.130000 196.760000 73.450000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 197.165000 73.450000 197.485000 ;
      LAYER met4 ;
        RECT 73.130000 197.165000 73.450000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 197.570000 73.450000 197.890000 ;
      LAYER met4 ;
        RECT 73.130000 197.570000 73.450000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 197.975000 73.450000 198.295000 ;
      LAYER met4 ;
        RECT 73.130000 197.975000 73.450000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 198.380000 73.450000 198.700000 ;
      LAYER met4 ;
        RECT 73.130000 198.380000 73.450000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 198.785000 73.450000 199.105000 ;
      LAYER met4 ;
        RECT 73.130000 198.785000 73.450000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 199.190000 73.450000 199.510000 ;
      LAYER met4 ;
        RECT 73.130000 199.190000 73.450000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 199.595000 73.450000 199.915000 ;
      LAYER met4 ;
        RECT 73.130000 199.595000 73.450000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 25.850000 73.450000 26.170000 ;
      LAYER met4 ;
        RECT 73.130000 25.850000 73.450000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 26.280000 73.450000 26.600000 ;
      LAYER met4 ;
        RECT 73.130000 26.280000 73.450000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 26.710000 73.450000 27.030000 ;
      LAYER met4 ;
        RECT 73.130000 26.710000 73.450000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 27.140000 73.450000 27.460000 ;
      LAYER met4 ;
        RECT 73.130000 27.140000 73.450000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 27.570000 73.450000 27.890000 ;
      LAYER met4 ;
        RECT 73.130000 27.570000 73.450000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 28.000000 73.450000 28.320000 ;
      LAYER met4 ;
        RECT 73.130000 28.000000 73.450000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 28.430000 73.450000 28.750000 ;
      LAYER met4 ;
        RECT 73.130000 28.430000 73.450000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 28.860000 73.450000 29.180000 ;
      LAYER met4 ;
        RECT 73.130000 28.860000 73.450000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 29.290000 73.450000 29.610000 ;
      LAYER met4 ;
        RECT 73.130000 29.290000 73.450000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 29.720000 73.450000 30.040000 ;
      LAYER met4 ;
        RECT 73.130000 29.720000 73.450000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 30.150000 73.450000 30.470000 ;
      LAYER met4 ;
        RECT 73.130000 30.150000 73.450000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 175.995000 73.390000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 176.395000 73.390000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 176.795000 73.390000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 177.195000 73.390000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 177.595000 73.390000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 177.995000 73.390000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 178.395000 73.390000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 178.795000 73.390000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 179.195000 73.390000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 179.595000 73.390000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 179.995000 73.390000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 180.395000 73.390000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 180.795000 73.390000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 181.195000 73.390000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 181.595000 73.390000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 181.995000 73.390000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 182.395000 73.390000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 182.795000 73.390000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 183.195000 73.390000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 183.595000 73.390000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 183.995000 73.390000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 184.395000 73.390000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 184.795000 73.390000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 185.195000 73.390000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 185.595000 73.390000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 185.995000 73.390000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 186.395000 73.390000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 186.795000 73.390000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 187.195000 73.390000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 187.595000 73.390000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 187.995000 73.390000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 188.395000 73.390000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 188.795000 73.390000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 189.195000 73.390000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 189.595000 73.390000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 189.995000 73.390000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 190.395000 73.390000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 190.795000 73.390000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 191.195000 73.390000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 191.595000 73.390000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 191.995000 73.390000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 192.395000 73.390000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 192.795000 73.390000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 193.195000 73.390000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 193.595000 73.390000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 193.995000 73.390000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 194.395000 73.390000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190000 194.795000 73.390000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 195.140000 73.850000 195.460000 ;
      LAYER met4 ;
        RECT 73.530000 195.140000 73.850000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 195.545000 73.850000 195.865000 ;
      LAYER met4 ;
        RECT 73.530000 195.545000 73.850000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 195.950000 73.850000 196.270000 ;
      LAYER met4 ;
        RECT 73.530000 195.950000 73.850000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 196.355000 73.850000 196.675000 ;
      LAYER met4 ;
        RECT 73.530000 196.355000 73.850000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 196.760000 73.850000 197.080000 ;
      LAYER met4 ;
        RECT 73.530000 196.760000 73.850000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 197.165000 73.850000 197.485000 ;
      LAYER met4 ;
        RECT 73.530000 197.165000 73.850000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 197.570000 73.850000 197.890000 ;
      LAYER met4 ;
        RECT 73.530000 197.570000 73.850000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 197.975000 73.850000 198.295000 ;
      LAYER met4 ;
        RECT 73.530000 197.975000 73.850000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 198.380000 73.850000 198.700000 ;
      LAYER met4 ;
        RECT 73.530000 198.380000 73.850000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 198.785000 73.850000 199.105000 ;
      LAYER met4 ;
        RECT 73.530000 198.785000 73.850000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 199.190000 73.850000 199.510000 ;
      LAYER met4 ;
        RECT 73.530000 199.190000 73.850000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 199.595000 73.850000 199.915000 ;
      LAYER met4 ;
        RECT 73.530000 199.595000 73.850000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 25.850000 73.855000 26.170000 ;
      LAYER met4 ;
        RECT 73.535000 25.850000 73.855000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 26.280000 73.855000 26.600000 ;
      LAYER met4 ;
        RECT 73.535000 26.280000 73.855000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 26.710000 73.855000 27.030000 ;
      LAYER met4 ;
        RECT 73.535000 26.710000 73.855000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 27.140000 73.855000 27.460000 ;
      LAYER met4 ;
        RECT 73.535000 27.140000 73.855000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 27.570000 73.855000 27.890000 ;
      LAYER met4 ;
        RECT 73.535000 27.570000 73.855000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 28.000000 73.855000 28.320000 ;
      LAYER met4 ;
        RECT 73.535000 28.000000 73.855000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 28.430000 73.855000 28.750000 ;
      LAYER met4 ;
        RECT 73.535000 28.430000 73.855000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 28.860000 73.855000 29.180000 ;
      LAYER met4 ;
        RECT 73.535000 28.860000 73.855000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 29.290000 73.855000 29.610000 ;
      LAYER met4 ;
        RECT 73.535000 29.290000 73.855000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 29.720000 73.855000 30.040000 ;
      LAYER met4 ;
        RECT 73.535000 29.720000 73.855000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 30.150000 73.855000 30.470000 ;
      LAYER met4 ;
        RECT 73.535000 30.150000 73.855000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 175.995000 73.790000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 176.395000 73.790000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 176.795000 73.790000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 177.195000 73.790000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 177.595000 73.790000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 177.995000 73.790000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 178.395000 73.790000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 178.795000 73.790000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 179.195000 73.790000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 179.595000 73.790000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 179.995000 73.790000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 180.395000 73.790000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 180.795000 73.790000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 181.195000 73.790000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 181.595000 73.790000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 181.995000 73.790000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 182.395000 73.790000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 182.795000 73.790000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 183.195000 73.790000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 183.595000 73.790000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 183.995000 73.790000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 184.395000 73.790000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 184.795000 73.790000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 185.195000 73.790000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 185.595000 73.790000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 185.995000 73.790000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 186.395000 73.790000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 186.795000 73.790000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 187.195000 73.790000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 187.595000 73.790000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 187.995000 73.790000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 188.395000 73.790000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 188.795000 73.790000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 189.195000 73.790000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 189.595000 73.790000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 189.995000 73.790000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 190.395000 73.790000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 190.795000 73.790000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 191.195000 73.790000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 191.595000 73.790000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 191.995000 73.790000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 192.395000 73.790000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 192.795000 73.790000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 193.195000 73.790000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 193.595000 73.790000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 193.995000 73.790000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 194.395000 73.790000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590000 194.795000 73.790000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 195.140000 74.250000 195.460000 ;
      LAYER met4 ;
        RECT 73.930000 195.140000 74.250000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 195.545000 74.250000 195.865000 ;
      LAYER met4 ;
        RECT 73.930000 195.545000 74.250000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 195.950000 74.250000 196.270000 ;
      LAYER met4 ;
        RECT 73.930000 195.950000 74.250000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 196.355000 74.250000 196.675000 ;
      LAYER met4 ;
        RECT 73.930000 196.355000 74.250000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 196.760000 74.250000 197.080000 ;
      LAYER met4 ;
        RECT 73.930000 196.760000 74.250000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 197.165000 74.250000 197.485000 ;
      LAYER met4 ;
        RECT 73.930000 197.165000 74.250000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 197.570000 74.250000 197.890000 ;
      LAYER met4 ;
        RECT 73.930000 197.570000 74.250000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 197.975000 74.250000 198.295000 ;
      LAYER met4 ;
        RECT 73.930000 197.975000 74.250000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 198.380000 74.250000 198.700000 ;
      LAYER met4 ;
        RECT 73.930000 198.380000 74.250000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 198.785000 74.250000 199.105000 ;
      LAYER met4 ;
        RECT 73.930000 198.785000 74.250000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 199.190000 74.250000 199.510000 ;
      LAYER met4 ;
        RECT 73.930000 199.190000 74.250000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930000 199.595000 74.250000 199.915000 ;
      LAYER met4 ;
        RECT 73.930000 199.595000 74.250000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 25.850000 74.260000 26.170000 ;
      LAYER met4 ;
        RECT 73.940000 25.850000 74.260000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 26.280000 74.260000 26.600000 ;
      LAYER met4 ;
        RECT 73.940000 26.280000 74.260000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 26.710000 74.260000 27.030000 ;
      LAYER met4 ;
        RECT 73.940000 26.710000 74.260000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 27.140000 74.260000 27.460000 ;
      LAYER met4 ;
        RECT 73.940000 27.140000 74.260000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 27.570000 74.260000 27.890000 ;
      LAYER met4 ;
        RECT 73.940000 27.570000 74.260000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 28.000000 74.260000 28.320000 ;
      LAYER met4 ;
        RECT 73.940000 28.000000 74.260000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 28.430000 74.260000 28.750000 ;
      LAYER met4 ;
        RECT 73.940000 28.430000 74.260000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 28.860000 74.260000 29.180000 ;
      LAYER met4 ;
        RECT 73.940000 28.860000 74.260000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 29.290000 74.260000 29.610000 ;
      LAYER met4 ;
        RECT 73.940000 29.290000 74.260000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 29.720000 74.260000 30.040000 ;
      LAYER met4 ;
        RECT 73.940000 29.720000 74.260000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 30.150000 74.260000 30.470000 ;
      LAYER met4 ;
        RECT 73.940000 30.150000 74.260000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 175.995000 74.190000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 176.395000 74.190000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 176.795000 74.190000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 177.195000 74.190000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 177.595000 74.190000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 177.995000 74.190000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 178.395000 74.190000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 178.795000 74.190000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 179.195000 74.190000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 179.595000 74.190000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 179.995000 74.190000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 180.395000 74.190000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 180.795000 74.190000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 181.195000 74.190000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 181.595000 74.190000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 181.995000 74.190000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 182.395000 74.190000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 182.795000 74.190000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 183.195000 74.190000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 183.595000 74.190000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 183.995000 74.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 184.395000 74.190000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 184.795000 74.190000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 185.195000 74.190000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 185.595000 74.190000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 185.995000 74.190000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 186.395000 74.190000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 186.795000 74.190000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 187.195000 74.190000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 187.595000 74.190000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 187.995000 74.190000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 188.395000 74.190000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 188.795000 74.190000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 189.195000 74.190000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 189.595000 74.190000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 189.995000 74.190000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 190.395000 74.190000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 190.795000 74.190000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 191.195000 74.190000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 191.595000 74.190000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 191.995000 74.190000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 192.395000 74.190000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 192.795000 74.190000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 193.195000 74.190000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 193.595000 74.190000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 193.995000 74.190000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.990000 194.395000 74.190000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 195.140000 8.545000 195.460000 ;
      LAYER met4 ;
        RECT 8.225000 195.140000 8.545000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 195.545000 8.545000 195.865000 ;
      LAYER met4 ;
        RECT 8.225000 195.545000 8.545000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 195.950000 8.545000 196.270000 ;
      LAYER met4 ;
        RECT 8.225000 195.950000 8.545000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 196.355000 8.545000 196.675000 ;
      LAYER met4 ;
        RECT 8.225000 196.355000 8.545000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 196.760000 8.545000 197.080000 ;
      LAYER met4 ;
        RECT 8.225000 196.760000 8.545000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 197.165000 8.545000 197.485000 ;
      LAYER met4 ;
        RECT 8.225000 197.165000 8.545000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 197.570000 8.545000 197.890000 ;
      LAYER met4 ;
        RECT 8.225000 197.570000 8.545000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 197.975000 8.545000 198.295000 ;
      LAYER met4 ;
        RECT 8.225000 197.975000 8.545000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 198.380000 8.545000 198.700000 ;
      LAYER met4 ;
        RECT 8.225000 198.380000 8.545000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 198.785000 8.545000 199.105000 ;
      LAYER met4 ;
        RECT 8.225000 198.785000 8.545000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 199.190000 8.545000 199.510000 ;
      LAYER met4 ;
        RECT 8.225000 199.190000 8.545000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225000 199.595000 8.545000 199.915000 ;
      LAYER met4 ;
        RECT 8.225000 199.595000 8.545000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 25.850000 8.570000 26.170000 ;
      LAYER met4 ;
        RECT 8.250000 25.850000 8.570000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 26.280000 8.570000 26.600000 ;
      LAYER met4 ;
        RECT 8.250000 26.280000 8.570000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 26.710000 8.570000 27.030000 ;
      LAYER met4 ;
        RECT 8.250000 26.710000 8.570000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 27.140000 8.570000 27.460000 ;
      LAYER met4 ;
        RECT 8.250000 27.140000 8.570000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 27.570000 8.570000 27.890000 ;
      LAYER met4 ;
        RECT 8.250000 27.570000 8.570000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 28.000000 8.570000 28.320000 ;
      LAYER met4 ;
        RECT 8.250000 28.000000 8.570000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 28.430000 8.570000 28.750000 ;
      LAYER met4 ;
        RECT 8.250000 28.430000 8.570000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 28.860000 8.570000 29.180000 ;
      LAYER met4 ;
        RECT 8.250000 28.860000 8.570000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 29.290000 8.570000 29.610000 ;
      LAYER met4 ;
        RECT 8.250000 29.290000 8.570000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 29.720000 8.570000 30.040000 ;
      LAYER met4 ;
        RECT 8.250000 29.720000 8.570000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 30.150000 8.570000 30.470000 ;
      LAYER met4 ;
        RECT 8.250000 30.150000 8.570000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 175.995000 8.485000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 176.395000 8.485000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 176.795000 8.485000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 177.195000 8.485000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 177.595000 8.485000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 177.995000 8.485000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 178.395000 8.485000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 178.795000 8.485000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 179.195000 8.485000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 179.595000 8.485000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 179.995000 8.485000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 180.395000 8.485000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 180.795000 8.485000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 181.195000 8.485000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 181.595000 8.485000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 181.995000 8.485000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 182.395000 8.485000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 182.795000 8.485000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 183.195000 8.485000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 183.595000 8.485000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 183.995000 8.485000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 184.395000 8.485000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 184.795000 8.485000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 185.195000 8.485000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 185.595000 8.485000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 185.995000 8.485000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 186.395000 8.485000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 186.795000 8.485000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 187.195000 8.485000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 187.595000 8.485000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 187.995000 8.485000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 188.395000 8.485000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 188.795000 8.485000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 189.195000 8.485000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 189.595000 8.485000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 189.995000 8.485000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 190.395000 8.485000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 190.795000 8.485000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 191.195000 8.485000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 191.595000 8.485000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 191.995000 8.485000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 192.395000 8.485000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 192.795000 8.485000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 193.195000 8.485000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 193.595000 8.485000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 193.995000 8.485000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 194.395000 8.485000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.285000 194.795000 8.485000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 195.140000 8.945000 195.460000 ;
      LAYER met4 ;
        RECT 8.625000 195.140000 8.945000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 195.545000 8.945000 195.865000 ;
      LAYER met4 ;
        RECT 8.625000 195.545000 8.945000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 195.950000 8.945000 196.270000 ;
      LAYER met4 ;
        RECT 8.625000 195.950000 8.945000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 196.355000 8.945000 196.675000 ;
      LAYER met4 ;
        RECT 8.625000 196.355000 8.945000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 196.760000 8.945000 197.080000 ;
      LAYER met4 ;
        RECT 8.625000 196.760000 8.945000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 197.165000 8.945000 197.485000 ;
      LAYER met4 ;
        RECT 8.625000 197.165000 8.945000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 197.570000 8.945000 197.890000 ;
      LAYER met4 ;
        RECT 8.625000 197.570000 8.945000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 197.975000 8.945000 198.295000 ;
      LAYER met4 ;
        RECT 8.625000 197.975000 8.945000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 198.380000 8.945000 198.700000 ;
      LAYER met4 ;
        RECT 8.625000 198.380000 8.945000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 198.785000 8.945000 199.105000 ;
      LAYER met4 ;
        RECT 8.625000 198.785000 8.945000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 199.190000 8.945000 199.510000 ;
      LAYER met4 ;
        RECT 8.625000 199.190000 8.945000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625000 199.595000 8.945000 199.915000 ;
      LAYER met4 ;
        RECT 8.625000 199.595000 8.945000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 25.850000 8.975000 26.170000 ;
      LAYER met4 ;
        RECT 8.655000 25.850000 8.975000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 26.280000 8.975000 26.600000 ;
      LAYER met4 ;
        RECT 8.655000 26.280000 8.975000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 26.710000 8.975000 27.030000 ;
      LAYER met4 ;
        RECT 8.655000 26.710000 8.975000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 27.140000 8.975000 27.460000 ;
      LAYER met4 ;
        RECT 8.655000 27.140000 8.975000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 27.570000 8.975000 27.890000 ;
      LAYER met4 ;
        RECT 8.655000 27.570000 8.975000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 28.000000 8.975000 28.320000 ;
      LAYER met4 ;
        RECT 8.655000 28.000000 8.975000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 28.430000 8.975000 28.750000 ;
      LAYER met4 ;
        RECT 8.655000 28.430000 8.975000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 28.860000 8.975000 29.180000 ;
      LAYER met4 ;
        RECT 8.655000 28.860000 8.975000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 29.290000 8.975000 29.610000 ;
      LAYER met4 ;
        RECT 8.655000 29.290000 8.975000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 29.720000 8.975000 30.040000 ;
      LAYER met4 ;
        RECT 8.655000 29.720000 8.975000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 30.150000 8.975000 30.470000 ;
      LAYER met4 ;
        RECT 8.655000 30.150000 8.975000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 175.995000 8.885000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 176.395000 8.885000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 176.795000 8.885000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 177.195000 8.885000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 177.595000 8.885000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 177.995000 8.885000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 178.395000 8.885000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 178.795000 8.885000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 179.195000 8.885000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 179.595000 8.885000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 179.995000 8.885000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 180.395000 8.885000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 180.795000 8.885000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 181.195000 8.885000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 181.595000 8.885000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 181.995000 8.885000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 182.395000 8.885000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 182.795000 8.885000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 183.195000 8.885000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 183.595000 8.885000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 183.995000 8.885000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 184.395000 8.885000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 184.795000 8.885000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 185.195000 8.885000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 185.595000 8.885000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 185.995000 8.885000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 186.395000 8.885000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 186.795000 8.885000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 187.195000 8.885000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 187.595000 8.885000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 187.995000 8.885000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 188.395000 8.885000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 188.795000 8.885000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 189.195000 8.885000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 189.595000 8.885000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 189.995000 8.885000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 190.395000 8.885000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 190.795000 8.885000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 191.195000 8.885000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 191.595000 8.885000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 191.995000 8.885000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 192.395000 8.885000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 192.795000 8.885000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 193.195000 8.885000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 193.595000 8.885000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 193.995000 8.885000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 194.395000 8.885000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.685000 194.795000 8.885000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 195.140000 9.345000 195.460000 ;
      LAYER met4 ;
        RECT 9.025000 195.140000 9.345000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 195.545000 9.345000 195.865000 ;
      LAYER met4 ;
        RECT 9.025000 195.545000 9.345000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 195.950000 9.345000 196.270000 ;
      LAYER met4 ;
        RECT 9.025000 195.950000 9.345000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 196.355000 9.345000 196.675000 ;
      LAYER met4 ;
        RECT 9.025000 196.355000 9.345000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 196.760000 9.345000 197.080000 ;
      LAYER met4 ;
        RECT 9.025000 196.760000 9.345000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 197.165000 9.345000 197.485000 ;
      LAYER met4 ;
        RECT 9.025000 197.165000 9.345000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 197.570000 9.345000 197.890000 ;
      LAYER met4 ;
        RECT 9.025000 197.570000 9.345000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 197.975000 9.345000 198.295000 ;
      LAYER met4 ;
        RECT 9.025000 197.975000 9.345000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 198.380000 9.345000 198.700000 ;
      LAYER met4 ;
        RECT 9.025000 198.380000 9.345000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 198.785000 9.345000 199.105000 ;
      LAYER met4 ;
        RECT 9.025000 198.785000 9.345000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 199.190000 9.345000 199.510000 ;
      LAYER met4 ;
        RECT 9.025000 199.190000 9.345000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025000 199.595000 9.345000 199.915000 ;
      LAYER met4 ;
        RECT 9.025000 199.595000 9.345000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 25.850000 9.380000 26.170000 ;
      LAYER met4 ;
        RECT 9.060000 25.850000 9.380000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 26.280000 9.380000 26.600000 ;
      LAYER met4 ;
        RECT 9.060000 26.280000 9.380000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 26.710000 9.380000 27.030000 ;
      LAYER met4 ;
        RECT 9.060000 26.710000 9.380000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 27.140000 9.380000 27.460000 ;
      LAYER met4 ;
        RECT 9.060000 27.140000 9.380000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 27.570000 9.380000 27.890000 ;
      LAYER met4 ;
        RECT 9.060000 27.570000 9.380000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 28.000000 9.380000 28.320000 ;
      LAYER met4 ;
        RECT 9.060000 28.000000 9.380000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 28.430000 9.380000 28.750000 ;
      LAYER met4 ;
        RECT 9.060000 28.430000 9.380000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 28.860000 9.380000 29.180000 ;
      LAYER met4 ;
        RECT 9.060000 28.860000 9.380000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 29.290000 9.380000 29.610000 ;
      LAYER met4 ;
        RECT 9.060000 29.290000 9.380000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 29.720000 9.380000 30.040000 ;
      LAYER met4 ;
        RECT 9.060000 29.720000 9.380000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 30.150000 9.380000 30.470000 ;
      LAYER met4 ;
        RECT 9.060000 30.150000 9.380000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 175.995000 9.285000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 176.395000 9.285000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 176.795000 9.285000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 177.195000 9.285000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 177.595000 9.285000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 177.995000 9.285000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 178.395000 9.285000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 178.795000 9.285000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 179.195000 9.285000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 179.595000 9.285000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 179.995000 9.285000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 180.395000 9.285000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 180.795000 9.285000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 181.195000 9.285000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 181.595000 9.285000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 181.995000 9.285000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 182.395000 9.285000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 182.795000 9.285000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 183.195000 9.285000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 183.595000 9.285000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 183.995000 9.285000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 184.395000 9.285000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 184.795000 9.285000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 185.195000 9.285000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 185.595000 9.285000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 185.995000 9.285000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 186.395000 9.285000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 186.795000 9.285000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 187.195000 9.285000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 187.595000 9.285000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 187.995000 9.285000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 188.395000 9.285000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 188.795000 9.285000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 189.195000 9.285000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 189.595000 9.285000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 189.995000 9.285000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 190.395000 9.285000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 190.795000 9.285000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 191.195000 9.285000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 191.595000 9.285000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 191.995000 9.285000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 192.395000 9.285000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 192.795000 9.285000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 193.195000 9.285000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 193.595000 9.285000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 193.995000 9.285000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 194.395000 9.285000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.085000 194.795000 9.285000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 195.140000 9.745000 195.460000 ;
      LAYER met4 ;
        RECT 9.425000 195.140000 9.745000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 195.545000 9.745000 195.865000 ;
      LAYER met4 ;
        RECT 9.425000 195.545000 9.745000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 195.950000 9.745000 196.270000 ;
      LAYER met4 ;
        RECT 9.425000 195.950000 9.745000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 196.355000 9.745000 196.675000 ;
      LAYER met4 ;
        RECT 9.425000 196.355000 9.745000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 196.760000 9.745000 197.080000 ;
      LAYER met4 ;
        RECT 9.425000 196.760000 9.745000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 197.165000 9.745000 197.485000 ;
      LAYER met4 ;
        RECT 9.425000 197.165000 9.745000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 197.570000 9.745000 197.890000 ;
      LAYER met4 ;
        RECT 9.425000 197.570000 9.745000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 197.975000 9.745000 198.295000 ;
      LAYER met4 ;
        RECT 9.425000 197.975000 9.745000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 198.380000 9.745000 198.700000 ;
      LAYER met4 ;
        RECT 9.425000 198.380000 9.745000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 198.785000 9.745000 199.105000 ;
      LAYER met4 ;
        RECT 9.425000 198.785000 9.745000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 199.190000 9.745000 199.510000 ;
      LAYER met4 ;
        RECT 9.425000 199.190000 9.745000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425000 199.595000 9.745000 199.915000 ;
      LAYER met4 ;
        RECT 9.425000 199.595000 9.745000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 25.850000 9.785000 26.170000 ;
      LAYER met4 ;
        RECT 9.465000 25.850000 9.785000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 26.280000 9.785000 26.600000 ;
      LAYER met4 ;
        RECT 9.465000 26.280000 9.785000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 26.710000 9.785000 27.030000 ;
      LAYER met4 ;
        RECT 9.465000 26.710000 9.785000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 27.140000 9.785000 27.460000 ;
      LAYER met4 ;
        RECT 9.465000 27.140000 9.785000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 27.570000 9.785000 27.890000 ;
      LAYER met4 ;
        RECT 9.465000 27.570000 9.785000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 28.000000 9.785000 28.320000 ;
      LAYER met4 ;
        RECT 9.465000 28.000000 9.785000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 28.430000 9.785000 28.750000 ;
      LAYER met4 ;
        RECT 9.465000 28.430000 9.785000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 28.860000 9.785000 29.180000 ;
      LAYER met4 ;
        RECT 9.465000 28.860000 9.785000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 29.290000 9.785000 29.610000 ;
      LAYER met4 ;
        RECT 9.465000 29.290000 9.785000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 29.720000 9.785000 30.040000 ;
      LAYER met4 ;
        RECT 9.465000 29.720000 9.785000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 30.150000 9.785000 30.470000 ;
      LAYER met4 ;
        RECT 9.465000 30.150000 9.785000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 175.995000 9.685000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 176.395000 9.685000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 176.795000 9.685000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 177.195000 9.685000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 177.595000 9.685000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 177.995000 9.685000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 178.395000 9.685000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 178.795000 9.685000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 179.195000 9.685000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 179.595000 9.685000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 179.995000 9.685000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 180.395000 9.685000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 180.795000 9.685000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 181.195000 9.685000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 181.595000 9.685000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 181.995000 9.685000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 182.395000 9.685000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 182.795000 9.685000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 183.195000 9.685000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 183.595000 9.685000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 183.995000 9.685000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 184.395000 9.685000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 184.795000 9.685000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 185.195000 9.685000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 185.595000 9.685000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 185.995000 9.685000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 186.395000 9.685000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 186.795000 9.685000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 187.195000 9.685000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 187.595000 9.685000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 187.995000 9.685000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 188.395000 9.685000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 188.795000 9.685000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 189.195000 9.685000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 189.595000 9.685000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 189.995000 9.685000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 190.395000 9.685000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 190.795000 9.685000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 191.195000 9.685000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 191.595000 9.685000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 191.995000 9.685000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 192.395000 9.685000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 192.795000 9.685000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 193.195000 9.685000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 193.595000 9.685000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 193.995000 9.685000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 194.395000 9.685000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.485000 194.795000 9.685000 194.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 195.140000 10.145000 195.460000 ;
      LAYER met4 ;
        RECT 9.825000 195.140000 10.145000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 195.545000 10.145000 195.865000 ;
      LAYER met4 ;
        RECT 9.825000 195.545000 10.145000 195.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 195.950000 10.145000 196.270000 ;
      LAYER met4 ;
        RECT 9.825000 195.950000 10.145000 196.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 196.355000 10.145000 196.675000 ;
      LAYER met4 ;
        RECT 9.825000 196.355000 10.145000 196.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 196.760000 10.145000 197.080000 ;
      LAYER met4 ;
        RECT 9.825000 196.760000 10.145000 197.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 197.165000 10.145000 197.485000 ;
      LAYER met4 ;
        RECT 9.825000 197.165000 10.145000 197.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 197.570000 10.145000 197.890000 ;
      LAYER met4 ;
        RECT 9.825000 197.570000 10.145000 197.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 197.975000 10.145000 198.295000 ;
      LAYER met4 ;
        RECT 9.825000 197.975000 10.145000 198.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 198.380000 10.145000 198.700000 ;
      LAYER met4 ;
        RECT 9.825000 198.380000 10.145000 198.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 198.785000 10.145000 199.105000 ;
      LAYER met4 ;
        RECT 9.825000 198.785000 10.145000 199.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 199.190000 10.145000 199.510000 ;
      LAYER met4 ;
        RECT 9.825000 199.190000 10.145000 199.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825000 199.595000 10.145000 199.915000 ;
      LAYER met4 ;
        RECT 9.825000 199.595000 10.145000 199.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 25.850000 10.190000 26.170000 ;
      LAYER met4 ;
        RECT 9.870000 25.850000 10.190000 26.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 26.280000 10.190000 26.600000 ;
      LAYER met4 ;
        RECT 9.870000 26.280000 10.190000 26.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 26.710000 10.190000 27.030000 ;
      LAYER met4 ;
        RECT 9.870000 26.710000 10.190000 27.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 27.140000 10.190000 27.460000 ;
      LAYER met4 ;
        RECT 9.870000 27.140000 10.190000 27.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 27.570000 10.190000 27.890000 ;
      LAYER met4 ;
        RECT 9.870000 27.570000 10.190000 27.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 28.000000 10.190000 28.320000 ;
      LAYER met4 ;
        RECT 9.870000 28.000000 10.190000 28.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 28.430000 10.190000 28.750000 ;
      LAYER met4 ;
        RECT 9.870000 28.430000 10.190000 28.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 28.860000 10.190000 29.180000 ;
      LAYER met4 ;
        RECT 9.870000 28.860000 10.190000 29.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 29.290000 10.190000 29.610000 ;
      LAYER met4 ;
        RECT 9.870000 29.290000 10.190000 29.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 29.720000 10.190000 30.040000 ;
      LAYER met4 ;
        RECT 9.870000 29.720000 10.190000 30.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 30.150000 10.190000 30.470000 ;
      LAYER met4 ;
        RECT 9.870000 30.150000 10.190000 30.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 175.995000 10.085000 176.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 176.395000 10.085000 176.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 176.795000 10.085000 176.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 177.195000 10.085000 177.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 177.595000 10.085000 177.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 177.995000 10.085000 178.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 178.395000 10.085000 178.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 178.795000 10.085000 178.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 179.195000 10.085000 179.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 179.595000 10.085000 179.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 179.995000 10.085000 180.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 180.395000 10.085000 180.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 180.795000 10.085000 180.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 181.195000 10.085000 181.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 181.595000 10.085000 181.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 181.995000 10.085000 182.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 182.395000 10.085000 182.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 182.795000 10.085000 182.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 183.195000 10.085000 183.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 183.595000 10.085000 183.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 183.995000 10.085000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 184.395000 10.085000 184.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 184.795000 10.085000 184.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 185.195000 10.085000 185.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 185.595000 10.085000 185.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 185.995000 10.085000 186.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 186.395000 10.085000 186.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 186.795000 10.085000 186.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 187.195000 10.085000 187.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 187.595000 10.085000 187.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 187.995000 10.085000 188.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 188.395000 10.085000 188.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 188.795000 10.085000 188.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 189.195000 10.085000 189.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 189.595000 10.085000 189.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 189.995000 10.085000 190.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 190.395000 10.085000 190.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 190.795000 10.085000 190.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 191.195000 10.085000 191.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 191.595000 10.085000 191.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 191.995000 10.085000 192.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 192.395000 10.085000 192.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 192.795000 10.085000 192.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 193.195000 10.085000 193.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 193.595000 10.085000 193.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 193.995000 10.085000 194.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 194.395000 10.085000 194.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.885000 194.795000 10.085000 194.995000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.525000 58.250000 0.845000 58.570000 ;
      LAYER met4 ;
        RECT 0.525000 58.250000 0.845000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 58.660000 0.845000 58.980000 ;
      LAYER met4 ;
        RECT 0.525000 58.660000 0.845000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 59.070000 0.845000 59.390000 ;
      LAYER met4 ;
        RECT 0.525000 59.070000 0.845000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 59.480000 0.845000 59.800000 ;
      LAYER met4 ;
        RECT 0.525000 59.480000 0.845000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 59.890000 0.845000 60.210000 ;
      LAYER met4 ;
        RECT 0.525000 59.890000 0.845000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 60.300000 0.845000 60.620000 ;
      LAYER met4 ;
        RECT 0.525000 60.300000 0.845000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 60.710000 0.845000 61.030000 ;
      LAYER met4 ;
        RECT 0.525000 60.710000 0.845000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 61.120000 0.845000 61.440000 ;
      LAYER met4 ;
        RECT 0.525000 61.120000 0.845000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 61.530000 0.845000 61.850000 ;
      LAYER met4 ;
        RECT 0.525000 61.530000 0.845000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 61.940000 0.845000 62.260000 ;
      LAYER met4 ;
        RECT 0.525000 61.940000 0.845000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 62.350000 0.845000 62.670000 ;
      LAYER met4 ;
        RECT 0.525000 62.350000 0.845000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 58.250000 1.255000 58.570000 ;
      LAYER met4 ;
        RECT 0.935000 58.250000 1.255000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 58.660000 1.255000 58.980000 ;
      LAYER met4 ;
        RECT 0.935000 58.660000 1.255000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 59.070000 1.255000 59.390000 ;
      LAYER met4 ;
        RECT 0.935000 59.070000 1.255000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 59.480000 1.255000 59.800000 ;
      LAYER met4 ;
        RECT 0.935000 59.480000 1.255000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 59.890000 1.255000 60.210000 ;
      LAYER met4 ;
        RECT 0.935000 59.890000 1.255000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 60.300000 1.255000 60.620000 ;
      LAYER met4 ;
        RECT 0.935000 60.300000 1.255000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 60.710000 1.255000 61.030000 ;
      LAYER met4 ;
        RECT 0.935000 60.710000 1.255000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 61.120000 1.255000 61.440000 ;
      LAYER met4 ;
        RECT 0.935000 61.120000 1.255000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 61.530000 1.255000 61.850000 ;
      LAYER met4 ;
        RECT 0.935000 61.530000 1.255000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 61.940000 1.255000 62.260000 ;
      LAYER met4 ;
        RECT 0.935000 61.940000 1.255000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 62.350000 1.255000 62.670000 ;
      LAYER met4 ;
        RECT 0.935000 62.350000 1.255000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 58.250000 1.665000 58.570000 ;
      LAYER met4 ;
        RECT 1.345000 58.250000 1.665000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 58.660000 1.665000 58.980000 ;
      LAYER met4 ;
        RECT 1.345000 58.660000 1.665000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 59.070000 1.665000 59.390000 ;
      LAYER met4 ;
        RECT 1.345000 59.070000 1.665000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 59.480000 1.665000 59.800000 ;
      LAYER met4 ;
        RECT 1.345000 59.480000 1.665000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 59.890000 1.665000 60.210000 ;
      LAYER met4 ;
        RECT 1.345000 59.890000 1.665000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 60.300000 1.665000 60.620000 ;
      LAYER met4 ;
        RECT 1.345000 60.300000 1.665000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 60.710000 1.665000 61.030000 ;
      LAYER met4 ;
        RECT 1.345000 60.710000 1.665000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 61.120000 1.665000 61.440000 ;
      LAYER met4 ;
        RECT 1.345000 61.120000 1.665000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 61.530000 1.665000 61.850000 ;
      LAYER met4 ;
        RECT 1.345000 61.530000 1.665000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 61.940000 1.665000 62.260000 ;
      LAYER met4 ;
        RECT 1.345000 61.940000 1.665000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 62.350000 1.665000 62.670000 ;
      LAYER met4 ;
        RECT 1.345000 62.350000 1.665000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 58.250000 2.075000 58.570000 ;
      LAYER met4 ;
        RECT 1.755000 58.250000 2.075000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 58.660000 2.075000 58.980000 ;
      LAYER met4 ;
        RECT 1.755000 58.660000 2.075000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 59.070000 2.075000 59.390000 ;
      LAYER met4 ;
        RECT 1.755000 59.070000 2.075000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 59.480000 2.075000 59.800000 ;
      LAYER met4 ;
        RECT 1.755000 59.480000 2.075000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 59.890000 2.075000 60.210000 ;
      LAYER met4 ;
        RECT 1.755000 59.890000 2.075000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 60.300000 2.075000 60.620000 ;
      LAYER met4 ;
        RECT 1.755000 60.300000 2.075000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 60.710000 2.075000 61.030000 ;
      LAYER met4 ;
        RECT 1.755000 60.710000 2.075000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 61.120000 2.075000 61.440000 ;
      LAYER met4 ;
        RECT 1.755000 61.120000 2.075000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 61.530000 2.075000 61.850000 ;
      LAYER met4 ;
        RECT 1.755000 61.530000 2.075000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 61.940000 2.075000 62.260000 ;
      LAYER met4 ;
        RECT 1.755000 61.940000 2.075000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 62.350000 2.075000 62.670000 ;
      LAYER met4 ;
        RECT 1.755000 62.350000 2.075000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 58.250000 10.595000 58.570000 ;
      LAYER met4 ;
        RECT 10.275000 58.250000 10.595000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 58.660000 10.595000 58.980000 ;
      LAYER met4 ;
        RECT 10.275000 58.660000 10.595000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 59.070000 10.595000 59.390000 ;
      LAYER met4 ;
        RECT 10.275000 59.070000 10.595000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 59.480000 10.595000 59.800000 ;
      LAYER met4 ;
        RECT 10.275000 59.480000 10.595000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 59.890000 10.595000 60.210000 ;
      LAYER met4 ;
        RECT 10.275000 59.890000 10.595000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 60.300000 10.595000 60.620000 ;
      LAYER met4 ;
        RECT 10.275000 60.300000 10.595000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 60.710000 10.595000 61.030000 ;
      LAYER met4 ;
        RECT 10.275000 60.710000 10.595000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 61.120000 10.595000 61.440000 ;
      LAYER met4 ;
        RECT 10.275000 61.120000 10.595000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 61.530000 10.595000 61.850000 ;
      LAYER met4 ;
        RECT 10.275000 61.530000 10.595000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 61.940000 10.595000 62.260000 ;
      LAYER met4 ;
        RECT 10.275000 61.940000 10.595000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 62.350000 10.595000 62.670000 ;
      LAYER met4 ;
        RECT 10.275000 62.350000 10.595000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 58.250000 11.000000 58.570000 ;
      LAYER met4 ;
        RECT 10.680000 58.250000 11.000000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 58.660000 11.000000 58.980000 ;
      LAYER met4 ;
        RECT 10.680000 58.660000 11.000000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 59.070000 11.000000 59.390000 ;
      LAYER met4 ;
        RECT 10.680000 59.070000 11.000000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 59.480000 11.000000 59.800000 ;
      LAYER met4 ;
        RECT 10.680000 59.480000 11.000000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 59.890000 11.000000 60.210000 ;
      LAYER met4 ;
        RECT 10.680000 59.890000 11.000000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 60.300000 11.000000 60.620000 ;
      LAYER met4 ;
        RECT 10.680000 60.300000 11.000000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 60.710000 11.000000 61.030000 ;
      LAYER met4 ;
        RECT 10.680000 60.710000 11.000000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 61.120000 11.000000 61.440000 ;
      LAYER met4 ;
        RECT 10.680000 61.120000 11.000000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 61.530000 11.000000 61.850000 ;
      LAYER met4 ;
        RECT 10.680000 61.530000 11.000000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 61.940000 11.000000 62.260000 ;
      LAYER met4 ;
        RECT 10.680000 61.940000 11.000000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 62.350000 11.000000 62.670000 ;
      LAYER met4 ;
        RECT 10.680000 62.350000 11.000000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 58.250000 11.405000 58.570000 ;
      LAYER met4 ;
        RECT 11.085000 58.250000 11.405000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 58.660000 11.405000 58.980000 ;
      LAYER met4 ;
        RECT 11.085000 58.660000 11.405000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 59.070000 11.405000 59.390000 ;
      LAYER met4 ;
        RECT 11.085000 59.070000 11.405000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 59.480000 11.405000 59.800000 ;
      LAYER met4 ;
        RECT 11.085000 59.480000 11.405000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 59.890000 11.405000 60.210000 ;
      LAYER met4 ;
        RECT 11.085000 59.890000 11.405000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 60.300000 11.405000 60.620000 ;
      LAYER met4 ;
        RECT 11.085000 60.300000 11.405000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 60.710000 11.405000 61.030000 ;
      LAYER met4 ;
        RECT 11.085000 60.710000 11.405000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 61.120000 11.405000 61.440000 ;
      LAYER met4 ;
        RECT 11.085000 61.120000 11.405000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 61.530000 11.405000 61.850000 ;
      LAYER met4 ;
        RECT 11.085000 61.530000 11.405000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 61.940000 11.405000 62.260000 ;
      LAYER met4 ;
        RECT 11.085000 61.940000 11.405000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 62.350000 11.405000 62.670000 ;
      LAYER met4 ;
        RECT 11.085000 62.350000 11.405000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 58.250000 11.810000 58.570000 ;
      LAYER met4 ;
        RECT 11.490000 58.250000 11.810000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 58.660000 11.810000 58.980000 ;
      LAYER met4 ;
        RECT 11.490000 58.660000 11.810000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 59.070000 11.810000 59.390000 ;
      LAYER met4 ;
        RECT 11.490000 59.070000 11.810000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 59.480000 11.810000 59.800000 ;
      LAYER met4 ;
        RECT 11.490000 59.480000 11.810000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 59.890000 11.810000 60.210000 ;
      LAYER met4 ;
        RECT 11.490000 59.890000 11.810000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 60.300000 11.810000 60.620000 ;
      LAYER met4 ;
        RECT 11.490000 60.300000 11.810000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 60.710000 11.810000 61.030000 ;
      LAYER met4 ;
        RECT 11.490000 60.710000 11.810000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 61.120000 11.810000 61.440000 ;
      LAYER met4 ;
        RECT 11.490000 61.120000 11.810000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 61.530000 11.810000 61.850000 ;
      LAYER met4 ;
        RECT 11.490000 61.530000 11.810000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 61.940000 11.810000 62.260000 ;
      LAYER met4 ;
        RECT 11.490000 61.940000 11.810000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 62.350000 11.810000 62.670000 ;
      LAYER met4 ;
        RECT 11.490000 62.350000 11.810000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 58.250000 12.215000 58.570000 ;
      LAYER met4 ;
        RECT 11.895000 58.250000 12.215000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 58.660000 12.215000 58.980000 ;
      LAYER met4 ;
        RECT 11.895000 58.660000 12.215000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 59.070000 12.215000 59.390000 ;
      LAYER met4 ;
        RECT 11.895000 59.070000 12.215000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 59.480000 12.215000 59.800000 ;
      LAYER met4 ;
        RECT 11.895000 59.480000 12.215000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 59.890000 12.215000 60.210000 ;
      LAYER met4 ;
        RECT 11.895000 59.890000 12.215000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 60.300000 12.215000 60.620000 ;
      LAYER met4 ;
        RECT 11.895000 60.300000 12.215000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 60.710000 12.215000 61.030000 ;
      LAYER met4 ;
        RECT 11.895000 60.710000 12.215000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 61.120000 12.215000 61.440000 ;
      LAYER met4 ;
        RECT 11.895000 61.120000 12.215000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 61.530000 12.215000 61.850000 ;
      LAYER met4 ;
        RECT 11.895000 61.530000 12.215000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 61.940000 12.215000 62.260000 ;
      LAYER met4 ;
        RECT 11.895000 61.940000 12.215000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 62.350000 12.215000 62.670000 ;
      LAYER met4 ;
        RECT 11.895000 62.350000 12.215000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 58.250000 12.620000 58.570000 ;
      LAYER met4 ;
        RECT 12.300000 58.250000 12.620000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 58.660000 12.620000 58.980000 ;
      LAYER met4 ;
        RECT 12.300000 58.660000 12.620000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 59.070000 12.620000 59.390000 ;
      LAYER met4 ;
        RECT 12.300000 59.070000 12.620000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 59.480000 12.620000 59.800000 ;
      LAYER met4 ;
        RECT 12.300000 59.480000 12.620000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 59.890000 12.620000 60.210000 ;
      LAYER met4 ;
        RECT 12.300000 59.890000 12.620000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 60.300000 12.620000 60.620000 ;
      LAYER met4 ;
        RECT 12.300000 60.300000 12.620000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 60.710000 12.620000 61.030000 ;
      LAYER met4 ;
        RECT 12.300000 60.710000 12.620000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 61.120000 12.620000 61.440000 ;
      LAYER met4 ;
        RECT 12.300000 61.120000 12.620000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 61.530000 12.620000 61.850000 ;
      LAYER met4 ;
        RECT 12.300000 61.530000 12.620000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 61.940000 12.620000 62.260000 ;
      LAYER met4 ;
        RECT 12.300000 61.940000 12.620000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 62.350000 12.620000 62.670000 ;
      LAYER met4 ;
        RECT 12.300000 62.350000 12.620000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 58.250000 13.025000 58.570000 ;
      LAYER met4 ;
        RECT 12.705000 58.250000 13.025000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 58.660000 13.025000 58.980000 ;
      LAYER met4 ;
        RECT 12.705000 58.660000 13.025000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 59.070000 13.025000 59.390000 ;
      LAYER met4 ;
        RECT 12.705000 59.070000 13.025000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 59.480000 13.025000 59.800000 ;
      LAYER met4 ;
        RECT 12.705000 59.480000 13.025000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 59.890000 13.025000 60.210000 ;
      LAYER met4 ;
        RECT 12.705000 59.890000 13.025000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 60.300000 13.025000 60.620000 ;
      LAYER met4 ;
        RECT 12.705000 60.300000 13.025000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 60.710000 13.025000 61.030000 ;
      LAYER met4 ;
        RECT 12.705000 60.710000 13.025000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 61.120000 13.025000 61.440000 ;
      LAYER met4 ;
        RECT 12.705000 61.120000 13.025000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 61.530000 13.025000 61.850000 ;
      LAYER met4 ;
        RECT 12.705000 61.530000 13.025000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 61.940000 13.025000 62.260000 ;
      LAYER met4 ;
        RECT 12.705000 61.940000 13.025000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 62.350000 13.025000 62.670000 ;
      LAYER met4 ;
        RECT 12.705000 62.350000 13.025000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 58.250000 13.430000 58.570000 ;
      LAYER met4 ;
        RECT 13.110000 58.250000 13.430000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 58.660000 13.430000 58.980000 ;
      LAYER met4 ;
        RECT 13.110000 58.660000 13.430000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 59.070000 13.430000 59.390000 ;
      LAYER met4 ;
        RECT 13.110000 59.070000 13.430000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 59.480000 13.430000 59.800000 ;
      LAYER met4 ;
        RECT 13.110000 59.480000 13.430000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 59.890000 13.430000 60.210000 ;
      LAYER met4 ;
        RECT 13.110000 59.890000 13.430000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 60.300000 13.430000 60.620000 ;
      LAYER met4 ;
        RECT 13.110000 60.300000 13.430000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 60.710000 13.430000 61.030000 ;
      LAYER met4 ;
        RECT 13.110000 60.710000 13.430000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 61.120000 13.430000 61.440000 ;
      LAYER met4 ;
        RECT 13.110000 61.120000 13.430000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 61.530000 13.430000 61.850000 ;
      LAYER met4 ;
        RECT 13.110000 61.530000 13.430000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 61.940000 13.430000 62.260000 ;
      LAYER met4 ;
        RECT 13.110000 61.940000 13.430000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 62.350000 13.430000 62.670000 ;
      LAYER met4 ;
        RECT 13.110000 62.350000 13.430000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 58.250000 13.835000 58.570000 ;
      LAYER met4 ;
        RECT 13.515000 58.250000 13.835000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 58.660000 13.835000 58.980000 ;
      LAYER met4 ;
        RECT 13.515000 58.660000 13.835000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 59.070000 13.835000 59.390000 ;
      LAYER met4 ;
        RECT 13.515000 59.070000 13.835000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 59.480000 13.835000 59.800000 ;
      LAYER met4 ;
        RECT 13.515000 59.480000 13.835000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 59.890000 13.835000 60.210000 ;
      LAYER met4 ;
        RECT 13.515000 59.890000 13.835000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 60.300000 13.835000 60.620000 ;
      LAYER met4 ;
        RECT 13.515000 60.300000 13.835000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 60.710000 13.835000 61.030000 ;
      LAYER met4 ;
        RECT 13.515000 60.710000 13.835000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 61.120000 13.835000 61.440000 ;
      LAYER met4 ;
        RECT 13.515000 61.120000 13.835000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 61.530000 13.835000 61.850000 ;
      LAYER met4 ;
        RECT 13.515000 61.530000 13.835000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 61.940000 13.835000 62.260000 ;
      LAYER met4 ;
        RECT 13.515000 61.940000 13.835000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 62.350000 13.835000 62.670000 ;
      LAYER met4 ;
        RECT 13.515000 62.350000 13.835000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 58.250000 14.240000 58.570000 ;
      LAYER met4 ;
        RECT 13.920000 58.250000 14.240000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 58.660000 14.240000 58.980000 ;
      LAYER met4 ;
        RECT 13.920000 58.660000 14.240000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 59.070000 14.240000 59.390000 ;
      LAYER met4 ;
        RECT 13.920000 59.070000 14.240000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 59.480000 14.240000 59.800000 ;
      LAYER met4 ;
        RECT 13.920000 59.480000 14.240000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 59.890000 14.240000 60.210000 ;
      LAYER met4 ;
        RECT 13.920000 59.890000 14.240000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 60.300000 14.240000 60.620000 ;
      LAYER met4 ;
        RECT 13.920000 60.300000 14.240000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 60.710000 14.240000 61.030000 ;
      LAYER met4 ;
        RECT 13.920000 60.710000 14.240000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 61.120000 14.240000 61.440000 ;
      LAYER met4 ;
        RECT 13.920000 61.120000 14.240000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 61.530000 14.240000 61.850000 ;
      LAYER met4 ;
        RECT 13.920000 61.530000 14.240000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 61.940000 14.240000 62.260000 ;
      LAYER met4 ;
        RECT 13.920000 61.940000 14.240000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 62.350000 14.240000 62.670000 ;
      LAYER met4 ;
        RECT 13.920000 62.350000 14.240000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 58.250000 14.645000 58.570000 ;
      LAYER met4 ;
        RECT 14.325000 58.250000 14.645000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 58.660000 14.645000 58.980000 ;
      LAYER met4 ;
        RECT 14.325000 58.660000 14.645000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 59.070000 14.645000 59.390000 ;
      LAYER met4 ;
        RECT 14.325000 59.070000 14.645000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 59.480000 14.645000 59.800000 ;
      LAYER met4 ;
        RECT 14.325000 59.480000 14.645000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 59.890000 14.645000 60.210000 ;
      LAYER met4 ;
        RECT 14.325000 59.890000 14.645000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 60.300000 14.645000 60.620000 ;
      LAYER met4 ;
        RECT 14.325000 60.300000 14.645000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 60.710000 14.645000 61.030000 ;
      LAYER met4 ;
        RECT 14.325000 60.710000 14.645000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 61.120000 14.645000 61.440000 ;
      LAYER met4 ;
        RECT 14.325000 61.120000 14.645000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 61.530000 14.645000 61.850000 ;
      LAYER met4 ;
        RECT 14.325000 61.530000 14.645000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 61.940000 14.645000 62.260000 ;
      LAYER met4 ;
        RECT 14.325000 61.940000 14.645000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 62.350000 14.645000 62.670000 ;
      LAYER met4 ;
        RECT 14.325000 62.350000 14.645000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 58.250000 15.050000 58.570000 ;
      LAYER met4 ;
        RECT 14.730000 58.250000 15.050000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 58.660000 15.050000 58.980000 ;
      LAYER met4 ;
        RECT 14.730000 58.660000 15.050000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 59.070000 15.050000 59.390000 ;
      LAYER met4 ;
        RECT 14.730000 59.070000 15.050000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 59.480000 15.050000 59.800000 ;
      LAYER met4 ;
        RECT 14.730000 59.480000 15.050000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 59.890000 15.050000 60.210000 ;
      LAYER met4 ;
        RECT 14.730000 59.890000 15.050000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 60.300000 15.050000 60.620000 ;
      LAYER met4 ;
        RECT 14.730000 60.300000 15.050000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 60.710000 15.050000 61.030000 ;
      LAYER met4 ;
        RECT 14.730000 60.710000 15.050000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 61.120000 15.050000 61.440000 ;
      LAYER met4 ;
        RECT 14.730000 61.120000 15.050000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 61.530000 15.050000 61.850000 ;
      LAYER met4 ;
        RECT 14.730000 61.530000 15.050000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 61.940000 15.050000 62.260000 ;
      LAYER met4 ;
        RECT 14.730000 61.940000 15.050000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 62.350000 15.050000 62.670000 ;
      LAYER met4 ;
        RECT 14.730000 62.350000 15.050000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 58.250000 15.455000 58.570000 ;
      LAYER met4 ;
        RECT 15.135000 58.250000 15.455000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 58.660000 15.455000 58.980000 ;
      LAYER met4 ;
        RECT 15.135000 58.660000 15.455000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 59.070000 15.455000 59.390000 ;
      LAYER met4 ;
        RECT 15.135000 59.070000 15.455000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 59.480000 15.455000 59.800000 ;
      LAYER met4 ;
        RECT 15.135000 59.480000 15.455000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 59.890000 15.455000 60.210000 ;
      LAYER met4 ;
        RECT 15.135000 59.890000 15.455000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 60.300000 15.455000 60.620000 ;
      LAYER met4 ;
        RECT 15.135000 60.300000 15.455000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 60.710000 15.455000 61.030000 ;
      LAYER met4 ;
        RECT 15.135000 60.710000 15.455000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 61.120000 15.455000 61.440000 ;
      LAYER met4 ;
        RECT 15.135000 61.120000 15.455000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 61.530000 15.455000 61.850000 ;
      LAYER met4 ;
        RECT 15.135000 61.530000 15.455000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 61.940000 15.455000 62.260000 ;
      LAYER met4 ;
        RECT 15.135000 61.940000 15.455000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 62.350000 15.455000 62.670000 ;
      LAYER met4 ;
        RECT 15.135000 62.350000 15.455000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 58.250000 15.860000 58.570000 ;
      LAYER met4 ;
        RECT 15.540000 58.250000 15.860000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 58.660000 15.860000 58.980000 ;
      LAYER met4 ;
        RECT 15.540000 58.660000 15.860000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 59.070000 15.860000 59.390000 ;
      LAYER met4 ;
        RECT 15.540000 59.070000 15.860000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 59.480000 15.860000 59.800000 ;
      LAYER met4 ;
        RECT 15.540000 59.480000 15.860000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 59.890000 15.860000 60.210000 ;
      LAYER met4 ;
        RECT 15.540000 59.890000 15.860000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 60.300000 15.860000 60.620000 ;
      LAYER met4 ;
        RECT 15.540000 60.300000 15.860000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 60.710000 15.860000 61.030000 ;
      LAYER met4 ;
        RECT 15.540000 60.710000 15.860000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 61.120000 15.860000 61.440000 ;
      LAYER met4 ;
        RECT 15.540000 61.120000 15.860000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 61.530000 15.860000 61.850000 ;
      LAYER met4 ;
        RECT 15.540000 61.530000 15.860000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 61.940000 15.860000 62.260000 ;
      LAYER met4 ;
        RECT 15.540000 61.940000 15.860000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 62.350000 15.860000 62.670000 ;
      LAYER met4 ;
        RECT 15.540000 62.350000 15.860000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 58.250000 16.265000 58.570000 ;
      LAYER met4 ;
        RECT 15.945000 58.250000 16.265000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 58.660000 16.265000 58.980000 ;
      LAYER met4 ;
        RECT 15.945000 58.660000 16.265000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 59.070000 16.265000 59.390000 ;
      LAYER met4 ;
        RECT 15.945000 59.070000 16.265000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 59.480000 16.265000 59.800000 ;
      LAYER met4 ;
        RECT 15.945000 59.480000 16.265000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 59.890000 16.265000 60.210000 ;
      LAYER met4 ;
        RECT 15.945000 59.890000 16.265000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 60.300000 16.265000 60.620000 ;
      LAYER met4 ;
        RECT 15.945000 60.300000 16.265000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 60.710000 16.265000 61.030000 ;
      LAYER met4 ;
        RECT 15.945000 60.710000 16.265000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 61.120000 16.265000 61.440000 ;
      LAYER met4 ;
        RECT 15.945000 61.120000 16.265000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 61.530000 16.265000 61.850000 ;
      LAYER met4 ;
        RECT 15.945000 61.530000 16.265000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 61.940000 16.265000 62.260000 ;
      LAYER met4 ;
        RECT 15.945000 61.940000 16.265000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 62.350000 16.265000 62.670000 ;
      LAYER met4 ;
        RECT 15.945000 62.350000 16.265000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 58.250000 16.670000 58.570000 ;
      LAYER met4 ;
        RECT 16.350000 58.250000 16.670000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 58.660000 16.670000 58.980000 ;
      LAYER met4 ;
        RECT 16.350000 58.660000 16.670000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 59.070000 16.670000 59.390000 ;
      LAYER met4 ;
        RECT 16.350000 59.070000 16.670000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 59.480000 16.670000 59.800000 ;
      LAYER met4 ;
        RECT 16.350000 59.480000 16.670000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 59.890000 16.670000 60.210000 ;
      LAYER met4 ;
        RECT 16.350000 59.890000 16.670000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 60.300000 16.670000 60.620000 ;
      LAYER met4 ;
        RECT 16.350000 60.300000 16.670000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 60.710000 16.670000 61.030000 ;
      LAYER met4 ;
        RECT 16.350000 60.710000 16.670000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 61.120000 16.670000 61.440000 ;
      LAYER met4 ;
        RECT 16.350000 61.120000 16.670000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 61.530000 16.670000 61.850000 ;
      LAYER met4 ;
        RECT 16.350000 61.530000 16.670000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 61.940000 16.670000 62.260000 ;
      LAYER met4 ;
        RECT 16.350000 61.940000 16.670000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 62.350000 16.670000 62.670000 ;
      LAYER met4 ;
        RECT 16.350000 62.350000 16.670000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 58.250000 17.075000 58.570000 ;
      LAYER met4 ;
        RECT 16.755000 58.250000 17.075000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 58.660000 17.075000 58.980000 ;
      LAYER met4 ;
        RECT 16.755000 58.660000 17.075000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 59.070000 17.075000 59.390000 ;
      LAYER met4 ;
        RECT 16.755000 59.070000 17.075000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 59.480000 17.075000 59.800000 ;
      LAYER met4 ;
        RECT 16.755000 59.480000 17.075000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 59.890000 17.075000 60.210000 ;
      LAYER met4 ;
        RECT 16.755000 59.890000 17.075000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 60.300000 17.075000 60.620000 ;
      LAYER met4 ;
        RECT 16.755000 60.300000 17.075000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 60.710000 17.075000 61.030000 ;
      LAYER met4 ;
        RECT 16.755000 60.710000 17.075000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 61.120000 17.075000 61.440000 ;
      LAYER met4 ;
        RECT 16.755000 61.120000 17.075000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 61.530000 17.075000 61.850000 ;
      LAYER met4 ;
        RECT 16.755000 61.530000 17.075000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 61.940000 17.075000 62.260000 ;
      LAYER met4 ;
        RECT 16.755000 61.940000 17.075000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 62.350000 17.075000 62.670000 ;
      LAYER met4 ;
        RECT 16.755000 62.350000 17.075000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 58.250000 17.480000 58.570000 ;
      LAYER met4 ;
        RECT 17.160000 58.250000 17.480000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 58.660000 17.480000 58.980000 ;
      LAYER met4 ;
        RECT 17.160000 58.660000 17.480000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 59.070000 17.480000 59.390000 ;
      LAYER met4 ;
        RECT 17.160000 59.070000 17.480000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 59.480000 17.480000 59.800000 ;
      LAYER met4 ;
        RECT 17.160000 59.480000 17.480000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 59.890000 17.480000 60.210000 ;
      LAYER met4 ;
        RECT 17.160000 59.890000 17.480000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 60.300000 17.480000 60.620000 ;
      LAYER met4 ;
        RECT 17.160000 60.300000 17.480000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 60.710000 17.480000 61.030000 ;
      LAYER met4 ;
        RECT 17.160000 60.710000 17.480000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 61.120000 17.480000 61.440000 ;
      LAYER met4 ;
        RECT 17.160000 61.120000 17.480000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 61.530000 17.480000 61.850000 ;
      LAYER met4 ;
        RECT 17.160000 61.530000 17.480000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 61.940000 17.480000 62.260000 ;
      LAYER met4 ;
        RECT 17.160000 61.940000 17.480000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 62.350000 17.480000 62.670000 ;
      LAYER met4 ;
        RECT 17.160000 62.350000 17.480000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 58.250000 17.885000 58.570000 ;
      LAYER met4 ;
        RECT 17.565000 58.250000 17.885000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 58.660000 17.885000 58.980000 ;
      LAYER met4 ;
        RECT 17.565000 58.660000 17.885000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 59.070000 17.885000 59.390000 ;
      LAYER met4 ;
        RECT 17.565000 59.070000 17.885000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 59.480000 17.885000 59.800000 ;
      LAYER met4 ;
        RECT 17.565000 59.480000 17.885000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 59.890000 17.885000 60.210000 ;
      LAYER met4 ;
        RECT 17.565000 59.890000 17.885000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 60.300000 17.885000 60.620000 ;
      LAYER met4 ;
        RECT 17.565000 60.300000 17.885000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 60.710000 17.885000 61.030000 ;
      LAYER met4 ;
        RECT 17.565000 60.710000 17.885000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 61.120000 17.885000 61.440000 ;
      LAYER met4 ;
        RECT 17.565000 61.120000 17.885000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 61.530000 17.885000 61.850000 ;
      LAYER met4 ;
        RECT 17.565000 61.530000 17.885000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 61.940000 17.885000 62.260000 ;
      LAYER met4 ;
        RECT 17.565000 61.940000 17.885000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 62.350000 17.885000 62.670000 ;
      LAYER met4 ;
        RECT 17.565000 62.350000 17.885000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 58.250000 18.290000 58.570000 ;
      LAYER met4 ;
        RECT 17.970000 58.250000 18.290000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 58.660000 18.290000 58.980000 ;
      LAYER met4 ;
        RECT 17.970000 58.660000 18.290000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 59.070000 18.290000 59.390000 ;
      LAYER met4 ;
        RECT 17.970000 59.070000 18.290000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 59.480000 18.290000 59.800000 ;
      LAYER met4 ;
        RECT 17.970000 59.480000 18.290000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 59.890000 18.290000 60.210000 ;
      LAYER met4 ;
        RECT 17.970000 59.890000 18.290000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 60.300000 18.290000 60.620000 ;
      LAYER met4 ;
        RECT 17.970000 60.300000 18.290000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 60.710000 18.290000 61.030000 ;
      LAYER met4 ;
        RECT 17.970000 60.710000 18.290000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 61.120000 18.290000 61.440000 ;
      LAYER met4 ;
        RECT 17.970000 61.120000 18.290000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 61.530000 18.290000 61.850000 ;
      LAYER met4 ;
        RECT 17.970000 61.530000 18.290000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 61.940000 18.290000 62.260000 ;
      LAYER met4 ;
        RECT 17.970000 61.940000 18.290000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 62.350000 18.290000 62.670000 ;
      LAYER met4 ;
        RECT 17.970000 62.350000 18.290000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 58.250000 18.695000 58.570000 ;
      LAYER met4 ;
        RECT 18.375000 58.250000 18.695000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 58.660000 18.695000 58.980000 ;
      LAYER met4 ;
        RECT 18.375000 58.660000 18.695000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 59.070000 18.695000 59.390000 ;
      LAYER met4 ;
        RECT 18.375000 59.070000 18.695000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 59.480000 18.695000 59.800000 ;
      LAYER met4 ;
        RECT 18.375000 59.480000 18.695000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 59.890000 18.695000 60.210000 ;
      LAYER met4 ;
        RECT 18.375000 59.890000 18.695000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 60.300000 18.695000 60.620000 ;
      LAYER met4 ;
        RECT 18.375000 60.300000 18.695000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 60.710000 18.695000 61.030000 ;
      LAYER met4 ;
        RECT 18.375000 60.710000 18.695000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 61.120000 18.695000 61.440000 ;
      LAYER met4 ;
        RECT 18.375000 61.120000 18.695000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 61.530000 18.695000 61.850000 ;
      LAYER met4 ;
        RECT 18.375000 61.530000 18.695000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 61.940000 18.695000 62.260000 ;
      LAYER met4 ;
        RECT 18.375000 61.940000 18.695000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 62.350000 18.695000 62.670000 ;
      LAYER met4 ;
        RECT 18.375000 62.350000 18.695000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 58.250000 19.100000 58.570000 ;
      LAYER met4 ;
        RECT 18.780000 58.250000 19.100000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 58.660000 19.100000 58.980000 ;
      LAYER met4 ;
        RECT 18.780000 58.660000 19.100000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 59.070000 19.100000 59.390000 ;
      LAYER met4 ;
        RECT 18.780000 59.070000 19.100000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 59.480000 19.100000 59.800000 ;
      LAYER met4 ;
        RECT 18.780000 59.480000 19.100000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 59.890000 19.100000 60.210000 ;
      LAYER met4 ;
        RECT 18.780000 59.890000 19.100000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 60.300000 19.100000 60.620000 ;
      LAYER met4 ;
        RECT 18.780000 60.300000 19.100000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 60.710000 19.100000 61.030000 ;
      LAYER met4 ;
        RECT 18.780000 60.710000 19.100000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 61.120000 19.100000 61.440000 ;
      LAYER met4 ;
        RECT 18.780000 61.120000 19.100000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 61.530000 19.100000 61.850000 ;
      LAYER met4 ;
        RECT 18.780000 61.530000 19.100000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 61.940000 19.100000 62.260000 ;
      LAYER met4 ;
        RECT 18.780000 61.940000 19.100000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 62.350000 19.100000 62.670000 ;
      LAYER met4 ;
        RECT 18.780000 62.350000 19.100000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 58.250000 19.505000 58.570000 ;
      LAYER met4 ;
        RECT 19.185000 58.250000 19.505000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 58.660000 19.505000 58.980000 ;
      LAYER met4 ;
        RECT 19.185000 58.660000 19.505000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 59.070000 19.505000 59.390000 ;
      LAYER met4 ;
        RECT 19.185000 59.070000 19.505000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 59.480000 19.505000 59.800000 ;
      LAYER met4 ;
        RECT 19.185000 59.480000 19.505000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 59.890000 19.505000 60.210000 ;
      LAYER met4 ;
        RECT 19.185000 59.890000 19.505000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 60.300000 19.505000 60.620000 ;
      LAYER met4 ;
        RECT 19.185000 60.300000 19.505000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 60.710000 19.505000 61.030000 ;
      LAYER met4 ;
        RECT 19.185000 60.710000 19.505000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 61.120000 19.505000 61.440000 ;
      LAYER met4 ;
        RECT 19.185000 61.120000 19.505000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 61.530000 19.505000 61.850000 ;
      LAYER met4 ;
        RECT 19.185000 61.530000 19.505000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 61.940000 19.505000 62.260000 ;
      LAYER met4 ;
        RECT 19.185000 61.940000 19.505000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 62.350000 19.505000 62.670000 ;
      LAYER met4 ;
        RECT 19.185000 62.350000 19.505000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 58.250000 19.910000 58.570000 ;
      LAYER met4 ;
        RECT 19.590000 58.250000 19.910000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 58.660000 19.910000 58.980000 ;
      LAYER met4 ;
        RECT 19.590000 58.660000 19.910000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 59.070000 19.910000 59.390000 ;
      LAYER met4 ;
        RECT 19.590000 59.070000 19.910000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 59.480000 19.910000 59.800000 ;
      LAYER met4 ;
        RECT 19.590000 59.480000 19.910000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 59.890000 19.910000 60.210000 ;
      LAYER met4 ;
        RECT 19.590000 59.890000 19.910000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 60.300000 19.910000 60.620000 ;
      LAYER met4 ;
        RECT 19.590000 60.300000 19.910000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 60.710000 19.910000 61.030000 ;
      LAYER met4 ;
        RECT 19.590000 60.710000 19.910000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 61.120000 19.910000 61.440000 ;
      LAYER met4 ;
        RECT 19.590000 61.120000 19.910000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 61.530000 19.910000 61.850000 ;
      LAYER met4 ;
        RECT 19.590000 61.530000 19.910000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 61.940000 19.910000 62.260000 ;
      LAYER met4 ;
        RECT 19.590000 61.940000 19.910000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 62.350000 19.910000 62.670000 ;
      LAYER met4 ;
        RECT 19.590000 62.350000 19.910000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 58.250000 20.315000 58.570000 ;
      LAYER met4 ;
        RECT 19.995000 58.250000 20.315000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 58.660000 20.315000 58.980000 ;
      LAYER met4 ;
        RECT 19.995000 58.660000 20.315000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 59.070000 20.315000 59.390000 ;
      LAYER met4 ;
        RECT 19.995000 59.070000 20.315000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 59.480000 20.315000 59.800000 ;
      LAYER met4 ;
        RECT 19.995000 59.480000 20.315000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 59.890000 20.315000 60.210000 ;
      LAYER met4 ;
        RECT 19.995000 59.890000 20.315000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 60.300000 20.315000 60.620000 ;
      LAYER met4 ;
        RECT 19.995000 60.300000 20.315000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 60.710000 20.315000 61.030000 ;
      LAYER met4 ;
        RECT 19.995000 60.710000 20.315000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 61.120000 20.315000 61.440000 ;
      LAYER met4 ;
        RECT 19.995000 61.120000 20.315000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 61.530000 20.315000 61.850000 ;
      LAYER met4 ;
        RECT 19.995000 61.530000 20.315000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 61.940000 20.315000 62.260000 ;
      LAYER met4 ;
        RECT 19.995000 61.940000 20.315000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 62.350000 20.315000 62.670000 ;
      LAYER met4 ;
        RECT 19.995000 62.350000 20.315000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 58.250000 2.485000 58.570000 ;
      LAYER met4 ;
        RECT 2.165000 58.250000 2.485000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 58.660000 2.485000 58.980000 ;
      LAYER met4 ;
        RECT 2.165000 58.660000 2.485000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 59.070000 2.485000 59.390000 ;
      LAYER met4 ;
        RECT 2.165000 59.070000 2.485000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 59.480000 2.485000 59.800000 ;
      LAYER met4 ;
        RECT 2.165000 59.480000 2.485000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 59.890000 2.485000 60.210000 ;
      LAYER met4 ;
        RECT 2.165000 59.890000 2.485000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 60.300000 2.485000 60.620000 ;
      LAYER met4 ;
        RECT 2.165000 60.300000 2.485000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 60.710000 2.485000 61.030000 ;
      LAYER met4 ;
        RECT 2.165000 60.710000 2.485000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 61.120000 2.485000 61.440000 ;
      LAYER met4 ;
        RECT 2.165000 61.120000 2.485000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 61.530000 2.485000 61.850000 ;
      LAYER met4 ;
        RECT 2.165000 61.530000 2.485000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 61.940000 2.485000 62.260000 ;
      LAYER met4 ;
        RECT 2.165000 61.940000 2.485000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 62.350000 2.485000 62.670000 ;
      LAYER met4 ;
        RECT 2.165000 62.350000 2.485000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 58.250000 2.895000 58.570000 ;
      LAYER met4 ;
        RECT 2.575000 58.250000 2.895000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 58.660000 2.895000 58.980000 ;
      LAYER met4 ;
        RECT 2.575000 58.660000 2.895000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 59.070000 2.895000 59.390000 ;
      LAYER met4 ;
        RECT 2.575000 59.070000 2.895000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 59.480000 2.895000 59.800000 ;
      LAYER met4 ;
        RECT 2.575000 59.480000 2.895000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 59.890000 2.895000 60.210000 ;
      LAYER met4 ;
        RECT 2.575000 59.890000 2.895000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 60.300000 2.895000 60.620000 ;
      LAYER met4 ;
        RECT 2.575000 60.300000 2.895000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 60.710000 2.895000 61.030000 ;
      LAYER met4 ;
        RECT 2.575000 60.710000 2.895000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 61.120000 2.895000 61.440000 ;
      LAYER met4 ;
        RECT 2.575000 61.120000 2.895000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 61.530000 2.895000 61.850000 ;
      LAYER met4 ;
        RECT 2.575000 61.530000 2.895000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 61.940000 2.895000 62.260000 ;
      LAYER met4 ;
        RECT 2.575000 61.940000 2.895000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 62.350000 2.895000 62.670000 ;
      LAYER met4 ;
        RECT 2.575000 62.350000 2.895000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 58.250000 3.305000 58.570000 ;
      LAYER met4 ;
        RECT 2.985000 58.250000 3.305000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 58.660000 3.305000 58.980000 ;
      LAYER met4 ;
        RECT 2.985000 58.660000 3.305000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 59.070000 3.305000 59.390000 ;
      LAYER met4 ;
        RECT 2.985000 59.070000 3.305000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 59.480000 3.305000 59.800000 ;
      LAYER met4 ;
        RECT 2.985000 59.480000 3.305000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 59.890000 3.305000 60.210000 ;
      LAYER met4 ;
        RECT 2.985000 59.890000 3.305000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 60.300000 3.305000 60.620000 ;
      LAYER met4 ;
        RECT 2.985000 60.300000 3.305000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 60.710000 3.305000 61.030000 ;
      LAYER met4 ;
        RECT 2.985000 60.710000 3.305000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 61.120000 3.305000 61.440000 ;
      LAYER met4 ;
        RECT 2.985000 61.120000 3.305000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 61.530000 3.305000 61.850000 ;
      LAYER met4 ;
        RECT 2.985000 61.530000 3.305000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 61.940000 3.305000 62.260000 ;
      LAYER met4 ;
        RECT 2.985000 61.940000 3.305000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 62.350000 3.305000 62.670000 ;
      LAYER met4 ;
        RECT 2.985000 62.350000 3.305000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 58.250000 20.720000 58.570000 ;
      LAYER met4 ;
        RECT 20.400000 58.250000 20.720000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 58.660000 20.720000 58.980000 ;
      LAYER met4 ;
        RECT 20.400000 58.660000 20.720000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 59.070000 20.720000 59.390000 ;
      LAYER met4 ;
        RECT 20.400000 59.070000 20.720000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 59.480000 20.720000 59.800000 ;
      LAYER met4 ;
        RECT 20.400000 59.480000 20.720000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 59.890000 20.720000 60.210000 ;
      LAYER met4 ;
        RECT 20.400000 59.890000 20.720000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 60.300000 20.720000 60.620000 ;
      LAYER met4 ;
        RECT 20.400000 60.300000 20.720000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 60.710000 20.720000 61.030000 ;
      LAYER met4 ;
        RECT 20.400000 60.710000 20.720000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 61.120000 20.720000 61.440000 ;
      LAYER met4 ;
        RECT 20.400000 61.120000 20.720000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 61.530000 20.720000 61.850000 ;
      LAYER met4 ;
        RECT 20.400000 61.530000 20.720000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 61.940000 20.720000 62.260000 ;
      LAYER met4 ;
        RECT 20.400000 61.940000 20.720000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 62.350000 20.720000 62.670000 ;
      LAYER met4 ;
        RECT 20.400000 62.350000 20.720000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 58.250000 21.125000 58.570000 ;
      LAYER met4 ;
        RECT 20.805000 58.250000 21.125000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 58.660000 21.125000 58.980000 ;
      LAYER met4 ;
        RECT 20.805000 58.660000 21.125000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 59.070000 21.125000 59.390000 ;
      LAYER met4 ;
        RECT 20.805000 59.070000 21.125000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 59.480000 21.125000 59.800000 ;
      LAYER met4 ;
        RECT 20.805000 59.480000 21.125000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 59.890000 21.125000 60.210000 ;
      LAYER met4 ;
        RECT 20.805000 59.890000 21.125000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 60.300000 21.125000 60.620000 ;
      LAYER met4 ;
        RECT 20.805000 60.300000 21.125000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 60.710000 21.125000 61.030000 ;
      LAYER met4 ;
        RECT 20.805000 60.710000 21.125000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 61.120000 21.125000 61.440000 ;
      LAYER met4 ;
        RECT 20.805000 61.120000 21.125000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 61.530000 21.125000 61.850000 ;
      LAYER met4 ;
        RECT 20.805000 61.530000 21.125000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 61.940000 21.125000 62.260000 ;
      LAYER met4 ;
        RECT 20.805000 61.940000 21.125000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 62.350000 21.125000 62.670000 ;
      LAYER met4 ;
        RECT 20.805000 62.350000 21.125000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 58.250000 21.530000 58.570000 ;
      LAYER met4 ;
        RECT 21.210000 58.250000 21.530000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 58.660000 21.530000 58.980000 ;
      LAYER met4 ;
        RECT 21.210000 58.660000 21.530000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 59.070000 21.530000 59.390000 ;
      LAYER met4 ;
        RECT 21.210000 59.070000 21.530000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 59.480000 21.530000 59.800000 ;
      LAYER met4 ;
        RECT 21.210000 59.480000 21.530000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 59.890000 21.530000 60.210000 ;
      LAYER met4 ;
        RECT 21.210000 59.890000 21.530000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 60.300000 21.530000 60.620000 ;
      LAYER met4 ;
        RECT 21.210000 60.300000 21.530000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 60.710000 21.530000 61.030000 ;
      LAYER met4 ;
        RECT 21.210000 60.710000 21.530000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 61.120000 21.530000 61.440000 ;
      LAYER met4 ;
        RECT 21.210000 61.120000 21.530000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 61.530000 21.530000 61.850000 ;
      LAYER met4 ;
        RECT 21.210000 61.530000 21.530000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 61.940000 21.530000 62.260000 ;
      LAYER met4 ;
        RECT 21.210000 61.940000 21.530000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 62.350000 21.530000 62.670000 ;
      LAYER met4 ;
        RECT 21.210000 62.350000 21.530000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 58.250000 21.935000 58.570000 ;
      LAYER met4 ;
        RECT 21.615000 58.250000 21.935000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 58.660000 21.935000 58.980000 ;
      LAYER met4 ;
        RECT 21.615000 58.660000 21.935000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 59.070000 21.935000 59.390000 ;
      LAYER met4 ;
        RECT 21.615000 59.070000 21.935000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 59.480000 21.935000 59.800000 ;
      LAYER met4 ;
        RECT 21.615000 59.480000 21.935000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 59.890000 21.935000 60.210000 ;
      LAYER met4 ;
        RECT 21.615000 59.890000 21.935000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 60.300000 21.935000 60.620000 ;
      LAYER met4 ;
        RECT 21.615000 60.300000 21.935000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 60.710000 21.935000 61.030000 ;
      LAYER met4 ;
        RECT 21.615000 60.710000 21.935000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 61.120000 21.935000 61.440000 ;
      LAYER met4 ;
        RECT 21.615000 61.120000 21.935000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 61.530000 21.935000 61.850000 ;
      LAYER met4 ;
        RECT 21.615000 61.530000 21.935000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 61.940000 21.935000 62.260000 ;
      LAYER met4 ;
        RECT 21.615000 61.940000 21.935000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 62.350000 21.935000 62.670000 ;
      LAYER met4 ;
        RECT 21.615000 62.350000 21.935000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 58.250000 22.340000 58.570000 ;
      LAYER met4 ;
        RECT 22.020000 58.250000 22.340000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 58.660000 22.340000 58.980000 ;
      LAYER met4 ;
        RECT 22.020000 58.660000 22.340000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 59.070000 22.340000 59.390000 ;
      LAYER met4 ;
        RECT 22.020000 59.070000 22.340000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 59.480000 22.340000 59.800000 ;
      LAYER met4 ;
        RECT 22.020000 59.480000 22.340000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 59.890000 22.340000 60.210000 ;
      LAYER met4 ;
        RECT 22.020000 59.890000 22.340000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 60.300000 22.340000 60.620000 ;
      LAYER met4 ;
        RECT 22.020000 60.300000 22.340000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 60.710000 22.340000 61.030000 ;
      LAYER met4 ;
        RECT 22.020000 60.710000 22.340000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 61.120000 22.340000 61.440000 ;
      LAYER met4 ;
        RECT 22.020000 61.120000 22.340000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 61.530000 22.340000 61.850000 ;
      LAYER met4 ;
        RECT 22.020000 61.530000 22.340000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 61.940000 22.340000 62.260000 ;
      LAYER met4 ;
        RECT 22.020000 61.940000 22.340000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 62.350000 22.340000 62.670000 ;
      LAYER met4 ;
        RECT 22.020000 62.350000 22.340000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 58.250000 22.745000 58.570000 ;
      LAYER met4 ;
        RECT 22.425000 58.250000 22.745000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 58.660000 22.745000 58.980000 ;
      LAYER met4 ;
        RECT 22.425000 58.660000 22.745000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 59.070000 22.745000 59.390000 ;
      LAYER met4 ;
        RECT 22.425000 59.070000 22.745000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 59.480000 22.745000 59.800000 ;
      LAYER met4 ;
        RECT 22.425000 59.480000 22.745000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 59.890000 22.745000 60.210000 ;
      LAYER met4 ;
        RECT 22.425000 59.890000 22.745000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 60.300000 22.745000 60.620000 ;
      LAYER met4 ;
        RECT 22.425000 60.300000 22.745000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 60.710000 22.745000 61.030000 ;
      LAYER met4 ;
        RECT 22.425000 60.710000 22.745000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 61.120000 22.745000 61.440000 ;
      LAYER met4 ;
        RECT 22.425000 61.120000 22.745000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 61.530000 22.745000 61.850000 ;
      LAYER met4 ;
        RECT 22.425000 61.530000 22.745000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 61.940000 22.745000 62.260000 ;
      LAYER met4 ;
        RECT 22.425000 61.940000 22.745000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 62.350000 22.745000 62.670000 ;
      LAYER met4 ;
        RECT 22.425000 62.350000 22.745000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 58.250000 23.150000 58.570000 ;
      LAYER met4 ;
        RECT 22.830000 58.250000 23.150000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 58.660000 23.150000 58.980000 ;
      LAYER met4 ;
        RECT 22.830000 58.660000 23.150000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 59.070000 23.150000 59.390000 ;
      LAYER met4 ;
        RECT 22.830000 59.070000 23.150000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 59.480000 23.150000 59.800000 ;
      LAYER met4 ;
        RECT 22.830000 59.480000 23.150000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 59.890000 23.150000 60.210000 ;
      LAYER met4 ;
        RECT 22.830000 59.890000 23.150000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 60.300000 23.150000 60.620000 ;
      LAYER met4 ;
        RECT 22.830000 60.300000 23.150000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 60.710000 23.150000 61.030000 ;
      LAYER met4 ;
        RECT 22.830000 60.710000 23.150000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 61.120000 23.150000 61.440000 ;
      LAYER met4 ;
        RECT 22.830000 61.120000 23.150000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 61.530000 23.150000 61.850000 ;
      LAYER met4 ;
        RECT 22.830000 61.530000 23.150000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 61.940000 23.150000 62.260000 ;
      LAYER met4 ;
        RECT 22.830000 61.940000 23.150000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 62.350000 23.150000 62.670000 ;
      LAYER met4 ;
        RECT 22.830000 62.350000 23.150000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 58.250000 23.555000 58.570000 ;
      LAYER met4 ;
        RECT 23.235000 58.250000 23.555000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 58.660000 23.555000 58.980000 ;
      LAYER met4 ;
        RECT 23.235000 58.660000 23.555000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 59.070000 23.555000 59.390000 ;
      LAYER met4 ;
        RECT 23.235000 59.070000 23.555000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 59.480000 23.555000 59.800000 ;
      LAYER met4 ;
        RECT 23.235000 59.480000 23.555000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 59.890000 23.555000 60.210000 ;
      LAYER met4 ;
        RECT 23.235000 59.890000 23.555000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 60.300000 23.555000 60.620000 ;
      LAYER met4 ;
        RECT 23.235000 60.300000 23.555000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 60.710000 23.555000 61.030000 ;
      LAYER met4 ;
        RECT 23.235000 60.710000 23.555000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 61.120000 23.555000 61.440000 ;
      LAYER met4 ;
        RECT 23.235000 61.120000 23.555000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 61.530000 23.555000 61.850000 ;
      LAYER met4 ;
        RECT 23.235000 61.530000 23.555000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 61.940000 23.555000 62.260000 ;
      LAYER met4 ;
        RECT 23.235000 61.940000 23.555000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 62.350000 23.555000 62.670000 ;
      LAYER met4 ;
        RECT 23.235000 62.350000 23.555000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 58.250000 23.960000 58.570000 ;
      LAYER met4 ;
        RECT 23.640000 58.250000 23.960000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 58.660000 23.960000 58.980000 ;
      LAYER met4 ;
        RECT 23.640000 58.660000 23.960000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 59.070000 23.960000 59.390000 ;
      LAYER met4 ;
        RECT 23.640000 59.070000 23.960000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 59.480000 23.960000 59.800000 ;
      LAYER met4 ;
        RECT 23.640000 59.480000 23.960000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 59.890000 23.960000 60.210000 ;
      LAYER met4 ;
        RECT 23.640000 59.890000 23.960000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 60.300000 23.960000 60.620000 ;
      LAYER met4 ;
        RECT 23.640000 60.300000 23.960000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 60.710000 23.960000 61.030000 ;
      LAYER met4 ;
        RECT 23.640000 60.710000 23.960000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 61.120000 23.960000 61.440000 ;
      LAYER met4 ;
        RECT 23.640000 61.120000 23.960000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 61.530000 23.960000 61.850000 ;
      LAYER met4 ;
        RECT 23.640000 61.530000 23.960000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 61.940000 23.960000 62.260000 ;
      LAYER met4 ;
        RECT 23.640000 61.940000 23.960000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 62.350000 23.960000 62.670000 ;
      LAYER met4 ;
        RECT 23.640000 62.350000 23.960000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 58.250000 24.365000 58.570000 ;
      LAYER met4 ;
        RECT 24.045000 58.250000 24.365000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 58.660000 24.365000 58.980000 ;
      LAYER met4 ;
        RECT 24.045000 58.660000 24.365000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 59.070000 24.365000 59.390000 ;
      LAYER met4 ;
        RECT 24.045000 59.070000 24.365000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 59.480000 24.365000 59.800000 ;
      LAYER met4 ;
        RECT 24.045000 59.480000 24.365000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 59.890000 24.365000 60.210000 ;
      LAYER met4 ;
        RECT 24.045000 59.890000 24.365000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 60.300000 24.365000 60.620000 ;
      LAYER met4 ;
        RECT 24.045000 60.300000 24.365000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 60.710000 24.365000 61.030000 ;
      LAYER met4 ;
        RECT 24.045000 60.710000 24.365000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 61.120000 24.365000 61.440000 ;
      LAYER met4 ;
        RECT 24.045000 61.120000 24.365000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 61.530000 24.365000 61.850000 ;
      LAYER met4 ;
        RECT 24.045000 61.530000 24.365000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 61.940000 24.365000 62.260000 ;
      LAYER met4 ;
        RECT 24.045000 61.940000 24.365000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 62.350000 24.365000 62.670000 ;
      LAYER met4 ;
        RECT 24.045000 62.350000 24.365000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 58.250000 3.710000 58.570000 ;
      LAYER met4 ;
        RECT 3.390000 58.250000 3.710000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 58.660000 3.710000 58.980000 ;
      LAYER met4 ;
        RECT 3.390000 58.660000 3.710000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 59.070000 3.710000 59.390000 ;
      LAYER met4 ;
        RECT 3.390000 59.070000 3.710000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 59.480000 3.710000 59.800000 ;
      LAYER met4 ;
        RECT 3.390000 59.480000 3.710000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 59.890000 3.710000 60.210000 ;
      LAYER met4 ;
        RECT 3.390000 59.890000 3.710000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 60.300000 3.710000 60.620000 ;
      LAYER met4 ;
        RECT 3.390000 60.300000 3.710000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 60.710000 3.710000 61.030000 ;
      LAYER met4 ;
        RECT 3.390000 60.710000 3.710000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 61.120000 3.710000 61.440000 ;
      LAYER met4 ;
        RECT 3.390000 61.120000 3.710000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 61.530000 3.710000 61.850000 ;
      LAYER met4 ;
        RECT 3.390000 61.530000 3.710000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 61.940000 3.710000 62.260000 ;
      LAYER met4 ;
        RECT 3.390000 61.940000 3.710000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 62.350000 3.710000 62.670000 ;
      LAYER met4 ;
        RECT 3.390000 62.350000 3.710000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 58.250000 4.115000 58.570000 ;
      LAYER met4 ;
        RECT 3.795000 58.250000 4.115000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 58.660000 4.115000 58.980000 ;
      LAYER met4 ;
        RECT 3.795000 58.660000 4.115000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 59.070000 4.115000 59.390000 ;
      LAYER met4 ;
        RECT 3.795000 59.070000 4.115000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 59.480000 4.115000 59.800000 ;
      LAYER met4 ;
        RECT 3.795000 59.480000 4.115000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 59.890000 4.115000 60.210000 ;
      LAYER met4 ;
        RECT 3.795000 59.890000 4.115000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 60.300000 4.115000 60.620000 ;
      LAYER met4 ;
        RECT 3.795000 60.300000 4.115000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 60.710000 4.115000 61.030000 ;
      LAYER met4 ;
        RECT 3.795000 60.710000 4.115000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 61.120000 4.115000 61.440000 ;
      LAYER met4 ;
        RECT 3.795000 61.120000 4.115000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 61.530000 4.115000 61.850000 ;
      LAYER met4 ;
        RECT 3.795000 61.530000 4.115000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 61.940000 4.115000 62.260000 ;
      LAYER met4 ;
        RECT 3.795000 61.940000 4.115000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 62.350000 4.115000 62.670000 ;
      LAYER met4 ;
        RECT 3.795000 62.350000 4.115000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 58.250000 4.520000 58.570000 ;
      LAYER met4 ;
        RECT 4.200000 58.250000 4.520000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 58.660000 4.520000 58.980000 ;
      LAYER met4 ;
        RECT 4.200000 58.660000 4.520000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 59.070000 4.520000 59.390000 ;
      LAYER met4 ;
        RECT 4.200000 59.070000 4.520000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 59.480000 4.520000 59.800000 ;
      LAYER met4 ;
        RECT 4.200000 59.480000 4.520000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 59.890000 4.520000 60.210000 ;
      LAYER met4 ;
        RECT 4.200000 59.890000 4.520000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 60.300000 4.520000 60.620000 ;
      LAYER met4 ;
        RECT 4.200000 60.300000 4.520000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 60.710000 4.520000 61.030000 ;
      LAYER met4 ;
        RECT 4.200000 60.710000 4.520000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 61.120000 4.520000 61.440000 ;
      LAYER met4 ;
        RECT 4.200000 61.120000 4.520000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 61.530000 4.520000 61.850000 ;
      LAYER met4 ;
        RECT 4.200000 61.530000 4.520000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 61.940000 4.520000 62.260000 ;
      LAYER met4 ;
        RECT 4.200000 61.940000 4.520000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 62.350000 4.520000 62.670000 ;
      LAYER met4 ;
        RECT 4.200000 62.350000 4.520000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 58.250000 4.925000 58.570000 ;
      LAYER met4 ;
        RECT 4.605000 58.250000 4.925000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 58.660000 4.925000 58.980000 ;
      LAYER met4 ;
        RECT 4.605000 58.660000 4.925000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 59.070000 4.925000 59.390000 ;
      LAYER met4 ;
        RECT 4.605000 59.070000 4.925000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 59.480000 4.925000 59.800000 ;
      LAYER met4 ;
        RECT 4.605000 59.480000 4.925000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 59.890000 4.925000 60.210000 ;
      LAYER met4 ;
        RECT 4.605000 59.890000 4.925000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 60.300000 4.925000 60.620000 ;
      LAYER met4 ;
        RECT 4.605000 60.300000 4.925000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 60.710000 4.925000 61.030000 ;
      LAYER met4 ;
        RECT 4.605000 60.710000 4.925000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 61.120000 4.925000 61.440000 ;
      LAYER met4 ;
        RECT 4.605000 61.120000 4.925000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 61.530000 4.925000 61.850000 ;
      LAYER met4 ;
        RECT 4.605000 61.530000 4.925000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 61.940000 4.925000 62.260000 ;
      LAYER met4 ;
        RECT 4.605000 61.940000 4.925000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 62.350000 4.925000 62.670000 ;
      LAYER met4 ;
        RECT 4.605000 62.350000 4.925000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 58.250000 5.330000 58.570000 ;
      LAYER met4 ;
        RECT 5.010000 58.250000 5.330000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 58.660000 5.330000 58.980000 ;
      LAYER met4 ;
        RECT 5.010000 58.660000 5.330000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 59.070000 5.330000 59.390000 ;
      LAYER met4 ;
        RECT 5.010000 59.070000 5.330000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 59.480000 5.330000 59.800000 ;
      LAYER met4 ;
        RECT 5.010000 59.480000 5.330000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 59.890000 5.330000 60.210000 ;
      LAYER met4 ;
        RECT 5.010000 59.890000 5.330000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 60.300000 5.330000 60.620000 ;
      LAYER met4 ;
        RECT 5.010000 60.300000 5.330000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 60.710000 5.330000 61.030000 ;
      LAYER met4 ;
        RECT 5.010000 60.710000 5.330000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 61.120000 5.330000 61.440000 ;
      LAYER met4 ;
        RECT 5.010000 61.120000 5.330000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 61.530000 5.330000 61.850000 ;
      LAYER met4 ;
        RECT 5.010000 61.530000 5.330000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 61.940000 5.330000 62.260000 ;
      LAYER met4 ;
        RECT 5.010000 61.940000 5.330000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 62.350000 5.330000 62.670000 ;
      LAYER met4 ;
        RECT 5.010000 62.350000 5.330000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 58.250000 5.735000 58.570000 ;
      LAYER met4 ;
        RECT 5.415000 58.250000 5.735000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 58.660000 5.735000 58.980000 ;
      LAYER met4 ;
        RECT 5.415000 58.660000 5.735000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 59.070000 5.735000 59.390000 ;
      LAYER met4 ;
        RECT 5.415000 59.070000 5.735000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 59.480000 5.735000 59.800000 ;
      LAYER met4 ;
        RECT 5.415000 59.480000 5.735000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 59.890000 5.735000 60.210000 ;
      LAYER met4 ;
        RECT 5.415000 59.890000 5.735000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 60.300000 5.735000 60.620000 ;
      LAYER met4 ;
        RECT 5.415000 60.300000 5.735000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 60.710000 5.735000 61.030000 ;
      LAYER met4 ;
        RECT 5.415000 60.710000 5.735000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 61.120000 5.735000 61.440000 ;
      LAYER met4 ;
        RECT 5.415000 61.120000 5.735000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 61.530000 5.735000 61.850000 ;
      LAYER met4 ;
        RECT 5.415000 61.530000 5.735000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 61.940000 5.735000 62.260000 ;
      LAYER met4 ;
        RECT 5.415000 61.940000 5.735000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 62.350000 5.735000 62.670000 ;
      LAYER met4 ;
        RECT 5.415000 62.350000 5.735000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 58.250000 6.140000 58.570000 ;
      LAYER met4 ;
        RECT 5.820000 58.250000 6.140000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 58.660000 6.140000 58.980000 ;
      LAYER met4 ;
        RECT 5.820000 58.660000 6.140000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 59.070000 6.140000 59.390000 ;
      LAYER met4 ;
        RECT 5.820000 59.070000 6.140000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 59.480000 6.140000 59.800000 ;
      LAYER met4 ;
        RECT 5.820000 59.480000 6.140000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 59.890000 6.140000 60.210000 ;
      LAYER met4 ;
        RECT 5.820000 59.890000 6.140000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 60.300000 6.140000 60.620000 ;
      LAYER met4 ;
        RECT 5.820000 60.300000 6.140000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 60.710000 6.140000 61.030000 ;
      LAYER met4 ;
        RECT 5.820000 60.710000 6.140000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 61.120000 6.140000 61.440000 ;
      LAYER met4 ;
        RECT 5.820000 61.120000 6.140000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 61.530000 6.140000 61.850000 ;
      LAYER met4 ;
        RECT 5.820000 61.530000 6.140000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 61.940000 6.140000 62.260000 ;
      LAYER met4 ;
        RECT 5.820000 61.940000 6.140000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 62.350000 6.140000 62.670000 ;
      LAYER met4 ;
        RECT 5.820000 62.350000 6.140000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 58.250000 50.740000 58.570000 ;
      LAYER met4 ;
        RECT 50.420000 58.250000 50.740000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 58.660000 50.740000 58.980000 ;
      LAYER met4 ;
        RECT 50.420000 58.660000 50.740000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 59.070000 50.740000 59.390000 ;
      LAYER met4 ;
        RECT 50.420000 59.070000 50.740000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 59.480000 50.740000 59.800000 ;
      LAYER met4 ;
        RECT 50.420000 59.480000 50.740000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 59.890000 50.740000 60.210000 ;
      LAYER met4 ;
        RECT 50.420000 59.890000 50.740000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 60.300000 50.740000 60.620000 ;
      LAYER met4 ;
        RECT 50.420000 60.300000 50.740000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 60.710000 50.740000 61.030000 ;
      LAYER met4 ;
        RECT 50.420000 60.710000 50.740000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 61.120000 50.740000 61.440000 ;
      LAYER met4 ;
        RECT 50.420000 61.120000 50.740000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 61.530000 50.740000 61.850000 ;
      LAYER met4 ;
        RECT 50.420000 61.530000 50.740000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 61.940000 50.740000 62.260000 ;
      LAYER met4 ;
        RECT 50.420000 61.940000 50.740000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 62.350000 50.740000 62.670000 ;
      LAYER met4 ;
        RECT 50.420000 62.350000 50.740000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 58.250000 51.150000 58.570000 ;
      LAYER met4 ;
        RECT 50.830000 58.250000 51.150000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 58.660000 51.150000 58.980000 ;
      LAYER met4 ;
        RECT 50.830000 58.660000 51.150000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 59.070000 51.150000 59.390000 ;
      LAYER met4 ;
        RECT 50.830000 59.070000 51.150000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 59.480000 51.150000 59.800000 ;
      LAYER met4 ;
        RECT 50.830000 59.480000 51.150000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 59.890000 51.150000 60.210000 ;
      LAYER met4 ;
        RECT 50.830000 59.890000 51.150000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 60.300000 51.150000 60.620000 ;
      LAYER met4 ;
        RECT 50.830000 60.300000 51.150000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 60.710000 51.150000 61.030000 ;
      LAYER met4 ;
        RECT 50.830000 60.710000 51.150000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 61.120000 51.150000 61.440000 ;
      LAYER met4 ;
        RECT 50.830000 61.120000 51.150000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 61.530000 51.150000 61.850000 ;
      LAYER met4 ;
        RECT 50.830000 61.530000 51.150000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 61.940000 51.150000 62.260000 ;
      LAYER met4 ;
        RECT 50.830000 61.940000 51.150000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 62.350000 51.150000 62.670000 ;
      LAYER met4 ;
        RECT 50.830000 62.350000 51.150000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 58.250000 51.560000 58.570000 ;
      LAYER met4 ;
        RECT 51.240000 58.250000 51.560000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 58.660000 51.560000 58.980000 ;
      LAYER met4 ;
        RECT 51.240000 58.660000 51.560000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 59.070000 51.560000 59.390000 ;
      LAYER met4 ;
        RECT 51.240000 59.070000 51.560000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 59.480000 51.560000 59.800000 ;
      LAYER met4 ;
        RECT 51.240000 59.480000 51.560000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 59.890000 51.560000 60.210000 ;
      LAYER met4 ;
        RECT 51.240000 59.890000 51.560000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 60.300000 51.560000 60.620000 ;
      LAYER met4 ;
        RECT 51.240000 60.300000 51.560000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 60.710000 51.560000 61.030000 ;
      LAYER met4 ;
        RECT 51.240000 60.710000 51.560000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 61.120000 51.560000 61.440000 ;
      LAYER met4 ;
        RECT 51.240000 61.120000 51.560000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 61.530000 51.560000 61.850000 ;
      LAYER met4 ;
        RECT 51.240000 61.530000 51.560000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 61.940000 51.560000 62.260000 ;
      LAYER met4 ;
        RECT 51.240000 61.940000 51.560000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 62.350000 51.560000 62.670000 ;
      LAYER met4 ;
        RECT 51.240000 62.350000 51.560000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 58.250000 51.970000 58.570000 ;
      LAYER met4 ;
        RECT 51.650000 58.250000 51.970000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 58.660000 51.970000 58.980000 ;
      LAYER met4 ;
        RECT 51.650000 58.660000 51.970000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 59.070000 51.970000 59.390000 ;
      LAYER met4 ;
        RECT 51.650000 59.070000 51.970000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 59.480000 51.970000 59.800000 ;
      LAYER met4 ;
        RECT 51.650000 59.480000 51.970000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 59.890000 51.970000 60.210000 ;
      LAYER met4 ;
        RECT 51.650000 59.890000 51.970000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 60.300000 51.970000 60.620000 ;
      LAYER met4 ;
        RECT 51.650000 60.300000 51.970000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 60.710000 51.970000 61.030000 ;
      LAYER met4 ;
        RECT 51.650000 60.710000 51.970000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 61.120000 51.970000 61.440000 ;
      LAYER met4 ;
        RECT 51.650000 61.120000 51.970000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 61.530000 51.970000 61.850000 ;
      LAYER met4 ;
        RECT 51.650000 61.530000 51.970000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 61.940000 51.970000 62.260000 ;
      LAYER met4 ;
        RECT 51.650000 61.940000 51.970000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 62.350000 51.970000 62.670000 ;
      LAYER met4 ;
        RECT 51.650000 62.350000 51.970000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 58.250000 52.380000 58.570000 ;
      LAYER met4 ;
        RECT 52.060000 58.250000 52.380000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 58.660000 52.380000 58.980000 ;
      LAYER met4 ;
        RECT 52.060000 58.660000 52.380000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 59.070000 52.380000 59.390000 ;
      LAYER met4 ;
        RECT 52.060000 59.070000 52.380000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 59.480000 52.380000 59.800000 ;
      LAYER met4 ;
        RECT 52.060000 59.480000 52.380000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 59.890000 52.380000 60.210000 ;
      LAYER met4 ;
        RECT 52.060000 59.890000 52.380000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 60.300000 52.380000 60.620000 ;
      LAYER met4 ;
        RECT 52.060000 60.300000 52.380000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 60.710000 52.380000 61.030000 ;
      LAYER met4 ;
        RECT 52.060000 60.710000 52.380000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 61.120000 52.380000 61.440000 ;
      LAYER met4 ;
        RECT 52.060000 61.120000 52.380000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 61.530000 52.380000 61.850000 ;
      LAYER met4 ;
        RECT 52.060000 61.530000 52.380000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 61.940000 52.380000 62.260000 ;
      LAYER met4 ;
        RECT 52.060000 61.940000 52.380000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 62.350000 52.380000 62.670000 ;
      LAYER met4 ;
        RECT 52.060000 62.350000 52.380000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 58.250000 52.790000 58.570000 ;
      LAYER met4 ;
        RECT 52.470000 58.250000 52.790000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 58.660000 52.790000 58.980000 ;
      LAYER met4 ;
        RECT 52.470000 58.660000 52.790000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 59.070000 52.790000 59.390000 ;
      LAYER met4 ;
        RECT 52.470000 59.070000 52.790000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 59.480000 52.790000 59.800000 ;
      LAYER met4 ;
        RECT 52.470000 59.480000 52.790000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 59.890000 52.790000 60.210000 ;
      LAYER met4 ;
        RECT 52.470000 59.890000 52.790000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 60.300000 52.790000 60.620000 ;
      LAYER met4 ;
        RECT 52.470000 60.300000 52.790000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 60.710000 52.790000 61.030000 ;
      LAYER met4 ;
        RECT 52.470000 60.710000 52.790000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 61.120000 52.790000 61.440000 ;
      LAYER met4 ;
        RECT 52.470000 61.120000 52.790000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 61.530000 52.790000 61.850000 ;
      LAYER met4 ;
        RECT 52.470000 61.530000 52.790000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 61.940000 52.790000 62.260000 ;
      LAYER met4 ;
        RECT 52.470000 61.940000 52.790000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 62.350000 52.790000 62.670000 ;
      LAYER met4 ;
        RECT 52.470000 62.350000 52.790000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 58.250000 53.200000 58.570000 ;
      LAYER met4 ;
        RECT 52.880000 58.250000 53.200000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 58.660000 53.200000 58.980000 ;
      LAYER met4 ;
        RECT 52.880000 58.660000 53.200000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 59.070000 53.200000 59.390000 ;
      LAYER met4 ;
        RECT 52.880000 59.070000 53.200000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 59.480000 53.200000 59.800000 ;
      LAYER met4 ;
        RECT 52.880000 59.480000 53.200000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 59.890000 53.200000 60.210000 ;
      LAYER met4 ;
        RECT 52.880000 59.890000 53.200000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 60.300000 53.200000 60.620000 ;
      LAYER met4 ;
        RECT 52.880000 60.300000 53.200000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 60.710000 53.200000 61.030000 ;
      LAYER met4 ;
        RECT 52.880000 60.710000 53.200000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 61.120000 53.200000 61.440000 ;
      LAYER met4 ;
        RECT 52.880000 61.120000 53.200000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 61.530000 53.200000 61.850000 ;
      LAYER met4 ;
        RECT 52.880000 61.530000 53.200000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 61.940000 53.200000 62.260000 ;
      LAYER met4 ;
        RECT 52.880000 61.940000 53.200000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 62.350000 53.200000 62.670000 ;
      LAYER met4 ;
        RECT 52.880000 62.350000 53.200000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 58.250000 53.605000 58.570000 ;
      LAYER met4 ;
        RECT 53.285000 58.250000 53.605000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 58.660000 53.605000 58.980000 ;
      LAYER met4 ;
        RECT 53.285000 58.660000 53.605000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 59.070000 53.605000 59.390000 ;
      LAYER met4 ;
        RECT 53.285000 59.070000 53.605000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 59.480000 53.605000 59.800000 ;
      LAYER met4 ;
        RECT 53.285000 59.480000 53.605000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 59.890000 53.605000 60.210000 ;
      LAYER met4 ;
        RECT 53.285000 59.890000 53.605000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 60.300000 53.605000 60.620000 ;
      LAYER met4 ;
        RECT 53.285000 60.300000 53.605000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 60.710000 53.605000 61.030000 ;
      LAYER met4 ;
        RECT 53.285000 60.710000 53.605000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 61.120000 53.605000 61.440000 ;
      LAYER met4 ;
        RECT 53.285000 61.120000 53.605000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 61.530000 53.605000 61.850000 ;
      LAYER met4 ;
        RECT 53.285000 61.530000 53.605000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 61.940000 53.605000 62.260000 ;
      LAYER met4 ;
        RECT 53.285000 61.940000 53.605000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 62.350000 53.605000 62.670000 ;
      LAYER met4 ;
        RECT 53.285000 62.350000 53.605000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 58.250000 54.010000 58.570000 ;
      LAYER met4 ;
        RECT 53.690000 58.250000 54.010000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 58.660000 54.010000 58.980000 ;
      LAYER met4 ;
        RECT 53.690000 58.660000 54.010000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 59.070000 54.010000 59.390000 ;
      LAYER met4 ;
        RECT 53.690000 59.070000 54.010000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 59.480000 54.010000 59.800000 ;
      LAYER met4 ;
        RECT 53.690000 59.480000 54.010000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 59.890000 54.010000 60.210000 ;
      LAYER met4 ;
        RECT 53.690000 59.890000 54.010000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 60.300000 54.010000 60.620000 ;
      LAYER met4 ;
        RECT 53.690000 60.300000 54.010000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 60.710000 54.010000 61.030000 ;
      LAYER met4 ;
        RECT 53.690000 60.710000 54.010000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 61.120000 54.010000 61.440000 ;
      LAYER met4 ;
        RECT 53.690000 61.120000 54.010000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 61.530000 54.010000 61.850000 ;
      LAYER met4 ;
        RECT 53.690000 61.530000 54.010000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 61.940000 54.010000 62.260000 ;
      LAYER met4 ;
        RECT 53.690000 61.940000 54.010000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 62.350000 54.010000 62.670000 ;
      LAYER met4 ;
        RECT 53.690000 62.350000 54.010000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 58.250000 54.415000 58.570000 ;
      LAYER met4 ;
        RECT 54.095000 58.250000 54.415000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 58.660000 54.415000 58.980000 ;
      LAYER met4 ;
        RECT 54.095000 58.660000 54.415000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 59.070000 54.415000 59.390000 ;
      LAYER met4 ;
        RECT 54.095000 59.070000 54.415000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 59.480000 54.415000 59.800000 ;
      LAYER met4 ;
        RECT 54.095000 59.480000 54.415000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 59.890000 54.415000 60.210000 ;
      LAYER met4 ;
        RECT 54.095000 59.890000 54.415000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 60.300000 54.415000 60.620000 ;
      LAYER met4 ;
        RECT 54.095000 60.300000 54.415000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 60.710000 54.415000 61.030000 ;
      LAYER met4 ;
        RECT 54.095000 60.710000 54.415000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 61.120000 54.415000 61.440000 ;
      LAYER met4 ;
        RECT 54.095000 61.120000 54.415000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 61.530000 54.415000 61.850000 ;
      LAYER met4 ;
        RECT 54.095000 61.530000 54.415000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 61.940000 54.415000 62.260000 ;
      LAYER met4 ;
        RECT 54.095000 61.940000 54.415000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 62.350000 54.415000 62.670000 ;
      LAYER met4 ;
        RECT 54.095000 62.350000 54.415000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 58.250000 54.820000 58.570000 ;
      LAYER met4 ;
        RECT 54.500000 58.250000 54.820000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 58.660000 54.820000 58.980000 ;
      LAYER met4 ;
        RECT 54.500000 58.660000 54.820000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 59.070000 54.820000 59.390000 ;
      LAYER met4 ;
        RECT 54.500000 59.070000 54.820000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 59.480000 54.820000 59.800000 ;
      LAYER met4 ;
        RECT 54.500000 59.480000 54.820000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 59.890000 54.820000 60.210000 ;
      LAYER met4 ;
        RECT 54.500000 59.890000 54.820000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 60.300000 54.820000 60.620000 ;
      LAYER met4 ;
        RECT 54.500000 60.300000 54.820000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 60.710000 54.820000 61.030000 ;
      LAYER met4 ;
        RECT 54.500000 60.710000 54.820000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 61.120000 54.820000 61.440000 ;
      LAYER met4 ;
        RECT 54.500000 61.120000 54.820000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 61.530000 54.820000 61.850000 ;
      LAYER met4 ;
        RECT 54.500000 61.530000 54.820000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 61.940000 54.820000 62.260000 ;
      LAYER met4 ;
        RECT 54.500000 61.940000 54.820000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 62.350000 54.820000 62.670000 ;
      LAYER met4 ;
        RECT 54.500000 62.350000 54.820000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 58.250000 55.225000 58.570000 ;
      LAYER met4 ;
        RECT 54.905000 58.250000 55.225000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 58.660000 55.225000 58.980000 ;
      LAYER met4 ;
        RECT 54.905000 58.660000 55.225000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 59.070000 55.225000 59.390000 ;
      LAYER met4 ;
        RECT 54.905000 59.070000 55.225000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 59.480000 55.225000 59.800000 ;
      LAYER met4 ;
        RECT 54.905000 59.480000 55.225000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 59.890000 55.225000 60.210000 ;
      LAYER met4 ;
        RECT 54.905000 59.890000 55.225000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 60.300000 55.225000 60.620000 ;
      LAYER met4 ;
        RECT 54.905000 60.300000 55.225000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 60.710000 55.225000 61.030000 ;
      LAYER met4 ;
        RECT 54.905000 60.710000 55.225000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 61.120000 55.225000 61.440000 ;
      LAYER met4 ;
        RECT 54.905000 61.120000 55.225000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 61.530000 55.225000 61.850000 ;
      LAYER met4 ;
        RECT 54.905000 61.530000 55.225000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 61.940000 55.225000 62.260000 ;
      LAYER met4 ;
        RECT 54.905000 61.940000 55.225000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 62.350000 55.225000 62.670000 ;
      LAYER met4 ;
        RECT 54.905000 62.350000 55.225000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 58.250000 55.630000 58.570000 ;
      LAYER met4 ;
        RECT 55.310000 58.250000 55.630000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 58.660000 55.630000 58.980000 ;
      LAYER met4 ;
        RECT 55.310000 58.660000 55.630000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 59.070000 55.630000 59.390000 ;
      LAYER met4 ;
        RECT 55.310000 59.070000 55.630000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 59.480000 55.630000 59.800000 ;
      LAYER met4 ;
        RECT 55.310000 59.480000 55.630000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 59.890000 55.630000 60.210000 ;
      LAYER met4 ;
        RECT 55.310000 59.890000 55.630000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 60.300000 55.630000 60.620000 ;
      LAYER met4 ;
        RECT 55.310000 60.300000 55.630000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 60.710000 55.630000 61.030000 ;
      LAYER met4 ;
        RECT 55.310000 60.710000 55.630000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 61.120000 55.630000 61.440000 ;
      LAYER met4 ;
        RECT 55.310000 61.120000 55.630000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 61.530000 55.630000 61.850000 ;
      LAYER met4 ;
        RECT 55.310000 61.530000 55.630000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 61.940000 55.630000 62.260000 ;
      LAYER met4 ;
        RECT 55.310000 61.940000 55.630000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 62.350000 55.630000 62.670000 ;
      LAYER met4 ;
        RECT 55.310000 62.350000 55.630000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 58.250000 56.035000 58.570000 ;
      LAYER met4 ;
        RECT 55.715000 58.250000 56.035000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 58.660000 56.035000 58.980000 ;
      LAYER met4 ;
        RECT 55.715000 58.660000 56.035000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 59.070000 56.035000 59.390000 ;
      LAYER met4 ;
        RECT 55.715000 59.070000 56.035000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 59.480000 56.035000 59.800000 ;
      LAYER met4 ;
        RECT 55.715000 59.480000 56.035000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 59.890000 56.035000 60.210000 ;
      LAYER met4 ;
        RECT 55.715000 59.890000 56.035000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 60.300000 56.035000 60.620000 ;
      LAYER met4 ;
        RECT 55.715000 60.300000 56.035000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 60.710000 56.035000 61.030000 ;
      LAYER met4 ;
        RECT 55.715000 60.710000 56.035000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 61.120000 56.035000 61.440000 ;
      LAYER met4 ;
        RECT 55.715000 61.120000 56.035000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 61.530000 56.035000 61.850000 ;
      LAYER met4 ;
        RECT 55.715000 61.530000 56.035000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 61.940000 56.035000 62.260000 ;
      LAYER met4 ;
        RECT 55.715000 61.940000 56.035000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 62.350000 56.035000 62.670000 ;
      LAYER met4 ;
        RECT 55.715000 62.350000 56.035000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 58.250000 56.440000 58.570000 ;
      LAYER met4 ;
        RECT 56.120000 58.250000 56.440000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 58.660000 56.440000 58.980000 ;
      LAYER met4 ;
        RECT 56.120000 58.660000 56.440000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 59.070000 56.440000 59.390000 ;
      LAYER met4 ;
        RECT 56.120000 59.070000 56.440000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 59.480000 56.440000 59.800000 ;
      LAYER met4 ;
        RECT 56.120000 59.480000 56.440000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 59.890000 56.440000 60.210000 ;
      LAYER met4 ;
        RECT 56.120000 59.890000 56.440000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 60.300000 56.440000 60.620000 ;
      LAYER met4 ;
        RECT 56.120000 60.300000 56.440000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 60.710000 56.440000 61.030000 ;
      LAYER met4 ;
        RECT 56.120000 60.710000 56.440000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 61.120000 56.440000 61.440000 ;
      LAYER met4 ;
        RECT 56.120000 61.120000 56.440000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 61.530000 56.440000 61.850000 ;
      LAYER met4 ;
        RECT 56.120000 61.530000 56.440000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 61.940000 56.440000 62.260000 ;
      LAYER met4 ;
        RECT 56.120000 61.940000 56.440000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 62.350000 56.440000 62.670000 ;
      LAYER met4 ;
        RECT 56.120000 62.350000 56.440000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 58.250000 56.845000 58.570000 ;
      LAYER met4 ;
        RECT 56.525000 58.250000 56.845000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 58.660000 56.845000 58.980000 ;
      LAYER met4 ;
        RECT 56.525000 58.660000 56.845000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 59.070000 56.845000 59.390000 ;
      LAYER met4 ;
        RECT 56.525000 59.070000 56.845000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 59.480000 56.845000 59.800000 ;
      LAYER met4 ;
        RECT 56.525000 59.480000 56.845000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 59.890000 56.845000 60.210000 ;
      LAYER met4 ;
        RECT 56.525000 59.890000 56.845000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 60.300000 56.845000 60.620000 ;
      LAYER met4 ;
        RECT 56.525000 60.300000 56.845000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 60.710000 56.845000 61.030000 ;
      LAYER met4 ;
        RECT 56.525000 60.710000 56.845000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 61.120000 56.845000 61.440000 ;
      LAYER met4 ;
        RECT 56.525000 61.120000 56.845000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 61.530000 56.845000 61.850000 ;
      LAYER met4 ;
        RECT 56.525000 61.530000 56.845000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 61.940000 56.845000 62.260000 ;
      LAYER met4 ;
        RECT 56.525000 61.940000 56.845000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 62.350000 56.845000 62.670000 ;
      LAYER met4 ;
        RECT 56.525000 62.350000 56.845000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 58.250000 57.250000 58.570000 ;
      LAYER met4 ;
        RECT 56.930000 58.250000 57.250000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 58.660000 57.250000 58.980000 ;
      LAYER met4 ;
        RECT 56.930000 58.660000 57.250000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 59.070000 57.250000 59.390000 ;
      LAYER met4 ;
        RECT 56.930000 59.070000 57.250000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 59.480000 57.250000 59.800000 ;
      LAYER met4 ;
        RECT 56.930000 59.480000 57.250000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 59.890000 57.250000 60.210000 ;
      LAYER met4 ;
        RECT 56.930000 59.890000 57.250000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 60.300000 57.250000 60.620000 ;
      LAYER met4 ;
        RECT 56.930000 60.300000 57.250000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 60.710000 57.250000 61.030000 ;
      LAYER met4 ;
        RECT 56.930000 60.710000 57.250000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 61.120000 57.250000 61.440000 ;
      LAYER met4 ;
        RECT 56.930000 61.120000 57.250000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 61.530000 57.250000 61.850000 ;
      LAYER met4 ;
        RECT 56.930000 61.530000 57.250000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 61.940000 57.250000 62.260000 ;
      LAYER met4 ;
        RECT 56.930000 61.940000 57.250000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 62.350000 57.250000 62.670000 ;
      LAYER met4 ;
        RECT 56.930000 62.350000 57.250000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 58.250000 57.655000 58.570000 ;
      LAYER met4 ;
        RECT 57.335000 58.250000 57.655000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 58.660000 57.655000 58.980000 ;
      LAYER met4 ;
        RECT 57.335000 58.660000 57.655000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 59.070000 57.655000 59.390000 ;
      LAYER met4 ;
        RECT 57.335000 59.070000 57.655000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 59.480000 57.655000 59.800000 ;
      LAYER met4 ;
        RECT 57.335000 59.480000 57.655000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 59.890000 57.655000 60.210000 ;
      LAYER met4 ;
        RECT 57.335000 59.890000 57.655000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 60.300000 57.655000 60.620000 ;
      LAYER met4 ;
        RECT 57.335000 60.300000 57.655000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 60.710000 57.655000 61.030000 ;
      LAYER met4 ;
        RECT 57.335000 60.710000 57.655000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 61.120000 57.655000 61.440000 ;
      LAYER met4 ;
        RECT 57.335000 61.120000 57.655000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 61.530000 57.655000 61.850000 ;
      LAYER met4 ;
        RECT 57.335000 61.530000 57.655000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 61.940000 57.655000 62.260000 ;
      LAYER met4 ;
        RECT 57.335000 61.940000 57.655000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 62.350000 57.655000 62.670000 ;
      LAYER met4 ;
        RECT 57.335000 62.350000 57.655000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 58.250000 58.060000 58.570000 ;
      LAYER met4 ;
        RECT 57.740000 58.250000 58.060000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 58.660000 58.060000 58.980000 ;
      LAYER met4 ;
        RECT 57.740000 58.660000 58.060000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 59.070000 58.060000 59.390000 ;
      LAYER met4 ;
        RECT 57.740000 59.070000 58.060000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 59.480000 58.060000 59.800000 ;
      LAYER met4 ;
        RECT 57.740000 59.480000 58.060000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 59.890000 58.060000 60.210000 ;
      LAYER met4 ;
        RECT 57.740000 59.890000 58.060000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 60.300000 58.060000 60.620000 ;
      LAYER met4 ;
        RECT 57.740000 60.300000 58.060000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 60.710000 58.060000 61.030000 ;
      LAYER met4 ;
        RECT 57.740000 60.710000 58.060000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 61.120000 58.060000 61.440000 ;
      LAYER met4 ;
        RECT 57.740000 61.120000 58.060000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 61.530000 58.060000 61.850000 ;
      LAYER met4 ;
        RECT 57.740000 61.530000 58.060000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 61.940000 58.060000 62.260000 ;
      LAYER met4 ;
        RECT 57.740000 61.940000 58.060000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 62.350000 58.060000 62.670000 ;
      LAYER met4 ;
        RECT 57.740000 62.350000 58.060000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 58.250000 58.465000 58.570000 ;
      LAYER met4 ;
        RECT 58.145000 58.250000 58.465000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 58.660000 58.465000 58.980000 ;
      LAYER met4 ;
        RECT 58.145000 58.660000 58.465000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 59.070000 58.465000 59.390000 ;
      LAYER met4 ;
        RECT 58.145000 59.070000 58.465000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 59.480000 58.465000 59.800000 ;
      LAYER met4 ;
        RECT 58.145000 59.480000 58.465000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 59.890000 58.465000 60.210000 ;
      LAYER met4 ;
        RECT 58.145000 59.890000 58.465000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 60.300000 58.465000 60.620000 ;
      LAYER met4 ;
        RECT 58.145000 60.300000 58.465000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 60.710000 58.465000 61.030000 ;
      LAYER met4 ;
        RECT 58.145000 60.710000 58.465000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 61.120000 58.465000 61.440000 ;
      LAYER met4 ;
        RECT 58.145000 61.120000 58.465000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 61.530000 58.465000 61.850000 ;
      LAYER met4 ;
        RECT 58.145000 61.530000 58.465000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 61.940000 58.465000 62.260000 ;
      LAYER met4 ;
        RECT 58.145000 61.940000 58.465000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 62.350000 58.465000 62.670000 ;
      LAYER met4 ;
        RECT 58.145000 62.350000 58.465000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 58.250000 58.870000 58.570000 ;
      LAYER met4 ;
        RECT 58.550000 58.250000 58.870000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 58.660000 58.870000 58.980000 ;
      LAYER met4 ;
        RECT 58.550000 58.660000 58.870000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 59.070000 58.870000 59.390000 ;
      LAYER met4 ;
        RECT 58.550000 59.070000 58.870000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 59.480000 58.870000 59.800000 ;
      LAYER met4 ;
        RECT 58.550000 59.480000 58.870000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 59.890000 58.870000 60.210000 ;
      LAYER met4 ;
        RECT 58.550000 59.890000 58.870000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 60.300000 58.870000 60.620000 ;
      LAYER met4 ;
        RECT 58.550000 60.300000 58.870000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 60.710000 58.870000 61.030000 ;
      LAYER met4 ;
        RECT 58.550000 60.710000 58.870000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 61.120000 58.870000 61.440000 ;
      LAYER met4 ;
        RECT 58.550000 61.120000 58.870000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 61.530000 58.870000 61.850000 ;
      LAYER met4 ;
        RECT 58.550000 61.530000 58.870000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 61.940000 58.870000 62.260000 ;
      LAYER met4 ;
        RECT 58.550000 61.940000 58.870000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 62.350000 58.870000 62.670000 ;
      LAYER met4 ;
        RECT 58.550000 62.350000 58.870000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 58.250000 59.275000 58.570000 ;
      LAYER met4 ;
        RECT 58.955000 58.250000 59.275000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 58.660000 59.275000 58.980000 ;
      LAYER met4 ;
        RECT 58.955000 58.660000 59.275000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 59.070000 59.275000 59.390000 ;
      LAYER met4 ;
        RECT 58.955000 59.070000 59.275000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 59.480000 59.275000 59.800000 ;
      LAYER met4 ;
        RECT 58.955000 59.480000 59.275000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 59.890000 59.275000 60.210000 ;
      LAYER met4 ;
        RECT 58.955000 59.890000 59.275000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 60.300000 59.275000 60.620000 ;
      LAYER met4 ;
        RECT 58.955000 60.300000 59.275000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 60.710000 59.275000 61.030000 ;
      LAYER met4 ;
        RECT 58.955000 60.710000 59.275000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 61.120000 59.275000 61.440000 ;
      LAYER met4 ;
        RECT 58.955000 61.120000 59.275000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 61.530000 59.275000 61.850000 ;
      LAYER met4 ;
        RECT 58.955000 61.530000 59.275000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 61.940000 59.275000 62.260000 ;
      LAYER met4 ;
        RECT 58.955000 61.940000 59.275000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 62.350000 59.275000 62.670000 ;
      LAYER met4 ;
        RECT 58.955000 62.350000 59.275000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 58.250000 59.680000 58.570000 ;
      LAYER met4 ;
        RECT 59.360000 58.250000 59.680000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 58.660000 59.680000 58.980000 ;
      LAYER met4 ;
        RECT 59.360000 58.660000 59.680000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 59.070000 59.680000 59.390000 ;
      LAYER met4 ;
        RECT 59.360000 59.070000 59.680000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 59.480000 59.680000 59.800000 ;
      LAYER met4 ;
        RECT 59.360000 59.480000 59.680000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 59.890000 59.680000 60.210000 ;
      LAYER met4 ;
        RECT 59.360000 59.890000 59.680000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 60.300000 59.680000 60.620000 ;
      LAYER met4 ;
        RECT 59.360000 60.300000 59.680000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 60.710000 59.680000 61.030000 ;
      LAYER met4 ;
        RECT 59.360000 60.710000 59.680000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 61.120000 59.680000 61.440000 ;
      LAYER met4 ;
        RECT 59.360000 61.120000 59.680000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 61.530000 59.680000 61.850000 ;
      LAYER met4 ;
        RECT 59.360000 61.530000 59.680000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 61.940000 59.680000 62.260000 ;
      LAYER met4 ;
        RECT 59.360000 61.940000 59.680000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 62.350000 59.680000 62.670000 ;
      LAYER met4 ;
        RECT 59.360000 62.350000 59.680000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 58.250000 60.085000 58.570000 ;
      LAYER met4 ;
        RECT 59.765000 58.250000 60.085000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 58.660000 60.085000 58.980000 ;
      LAYER met4 ;
        RECT 59.765000 58.660000 60.085000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 59.070000 60.085000 59.390000 ;
      LAYER met4 ;
        RECT 59.765000 59.070000 60.085000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 59.480000 60.085000 59.800000 ;
      LAYER met4 ;
        RECT 59.765000 59.480000 60.085000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 59.890000 60.085000 60.210000 ;
      LAYER met4 ;
        RECT 59.765000 59.890000 60.085000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 60.300000 60.085000 60.620000 ;
      LAYER met4 ;
        RECT 59.765000 60.300000 60.085000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 60.710000 60.085000 61.030000 ;
      LAYER met4 ;
        RECT 59.765000 60.710000 60.085000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 61.120000 60.085000 61.440000 ;
      LAYER met4 ;
        RECT 59.765000 61.120000 60.085000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 61.530000 60.085000 61.850000 ;
      LAYER met4 ;
        RECT 59.765000 61.530000 60.085000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 61.940000 60.085000 62.260000 ;
      LAYER met4 ;
        RECT 59.765000 61.940000 60.085000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 62.350000 60.085000 62.670000 ;
      LAYER met4 ;
        RECT 59.765000 62.350000 60.085000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 58.250000 6.545000 58.570000 ;
      LAYER met4 ;
        RECT 6.225000 58.250000 6.545000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 58.660000 6.545000 58.980000 ;
      LAYER met4 ;
        RECT 6.225000 58.660000 6.545000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 59.070000 6.545000 59.390000 ;
      LAYER met4 ;
        RECT 6.225000 59.070000 6.545000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 59.480000 6.545000 59.800000 ;
      LAYER met4 ;
        RECT 6.225000 59.480000 6.545000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 59.890000 6.545000 60.210000 ;
      LAYER met4 ;
        RECT 6.225000 59.890000 6.545000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 60.300000 6.545000 60.620000 ;
      LAYER met4 ;
        RECT 6.225000 60.300000 6.545000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 60.710000 6.545000 61.030000 ;
      LAYER met4 ;
        RECT 6.225000 60.710000 6.545000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 61.120000 6.545000 61.440000 ;
      LAYER met4 ;
        RECT 6.225000 61.120000 6.545000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 61.530000 6.545000 61.850000 ;
      LAYER met4 ;
        RECT 6.225000 61.530000 6.545000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 61.940000 6.545000 62.260000 ;
      LAYER met4 ;
        RECT 6.225000 61.940000 6.545000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 62.350000 6.545000 62.670000 ;
      LAYER met4 ;
        RECT 6.225000 62.350000 6.545000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 58.250000 6.950000 58.570000 ;
      LAYER met4 ;
        RECT 6.630000 58.250000 6.950000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 58.660000 6.950000 58.980000 ;
      LAYER met4 ;
        RECT 6.630000 58.660000 6.950000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 59.070000 6.950000 59.390000 ;
      LAYER met4 ;
        RECT 6.630000 59.070000 6.950000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 59.480000 6.950000 59.800000 ;
      LAYER met4 ;
        RECT 6.630000 59.480000 6.950000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 59.890000 6.950000 60.210000 ;
      LAYER met4 ;
        RECT 6.630000 59.890000 6.950000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 60.300000 6.950000 60.620000 ;
      LAYER met4 ;
        RECT 6.630000 60.300000 6.950000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 60.710000 6.950000 61.030000 ;
      LAYER met4 ;
        RECT 6.630000 60.710000 6.950000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 61.120000 6.950000 61.440000 ;
      LAYER met4 ;
        RECT 6.630000 61.120000 6.950000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 61.530000 6.950000 61.850000 ;
      LAYER met4 ;
        RECT 6.630000 61.530000 6.950000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 61.940000 6.950000 62.260000 ;
      LAYER met4 ;
        RECT 6.630000 61.940000 6.950000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 62.350000 6.950000 62.670000 ;
      LAYER met4 ;
        RECT 6.630000 62.350000 6.950000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 58.250000 60.490000 58.570000 ;
      LAYER met4 ;
        RECT 60.170000 58.250000 60.490000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 58.660000 60.490000 58.980000 ;
      LAYER met4 ;
        RECT 60.170000 58.660000 60.490000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 59.070000 60.490000 59.390000 ;
      LAYER met4 ;
        RECT 60.170000 59.070000 60.490000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 59.480000 60.490000 59.800000 ;
      LAYER met4 ;
        RECT 60.170000 59.480000 60.490000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 59.890000 60.490000 60.210000 ;
      LAYER met4 ;
        RECT 60.170000 59.890000 60.490000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 60.300000 60.490000 60.620000 ;
      LAYER met4 ;
        RECT 60.170000 60.300000 60.490000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 60.710000 60.490000 61.030000 ;
      LAYER met4 ;
        RECT 60.170000 60.710000 60.490000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 61.120000 60.490000 61.440000 ;
      LAYER met4 ;
        RECT 60.170000 61.120000 60.490000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 61.530000 60.490000 61.850000 ;
      LAYER met4 ;
        RECT 60.170000 61.530000 60.490000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 61.940000 60.490000 62.260000 ;
      LAYER met4 ;
        RECT 60.170000 61.940000 60.490000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 62.350000 60.490000 62.670000 ;
      LAYER met4 ;
        RECT 60.170000 62.350000 60.490000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 58.250000 60.895000 58.570000 ;
      LAYER met4 ;
        RECT 60.575000 58.250000 60.895000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 58.660000 60.895000 58.980000 ;
      LAYER met4 ;
        RECT 60.575000 58.660000 60.895000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 59.070000 60.895000 59.390000 ;
      LAYER met4 ;
        RECT 60.575000 59.070000 60.895000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 59.480000 60.895000 59.800000 ;
      LAYER met4 ;
        RECT 60.575000 59.480000 60.895000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 59.890000 60.895000 60.210000 ;
      LAYER met4 ;
        RECT 60.575000 59.890000 60.895000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 60.300000 60.895000 60.620000 ;
      LAYER met4 ;
        RECT 60.575000 60.300000 60.895000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 60.710000 60.895000 61.030000 ;
      LAYER met4 ;
        RECT 60.575000 60.710000 60.895000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 61.120000 60.895000 61.440000 ;
      LAYER met4 ;
        RECT 60.575000 61.120000 60.895000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 61.530000 60.895000 61.850000 ;
      LAYER met4 ;
        RECT 60.575000 61.530000 60.895000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 61.940000 60.895000 62.260000 ;
      LAYER met4 ;
        RECT 60.575000 61.940000 60.895000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 62.350000 60.895000 62.670000 ;
      LAYER met4 ;
        RECT 60.575000 62.350000 60.895000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 58.250000 61.300000 58.570000 ;
      LAYER met4 ;
        RECT 60.980000 58.250000 61.300000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 58.660000 61.300000 58.980000 ;
      LAYER met4 ;
        RECT 60.980000 58.660000 61.300000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 59.070000 61.300000 59.390000 ;
      LAYER met4 ;
        RECT 60.980000 59.070000 61.300000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 59.480000 61.300000 59.800000 ;
      LAYER met4 ;
        RECT 60.980000 59.480000 61.300000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 59.890000 61.300000 60.210000 ;
      LAYER met4 ;
        RECT 60.980000 59.890000 61.300000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 60.300000 61.300000 60.620000 ;
      LAYER met4 ;
        RECT 60.980000 60.300000 61.300000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 60.710000 61.300000 61.030000 ;
      LAYER met4 ;
        RECT 60.980000 60.710000 61.300000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 61.120000 61.300000 61.440000 ;
      LAYER met4 ;
        RECT 60.980000 61.120000 61.300000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 61.530000 61.300000 61.850000 ;
      LAYER met4 ;
        RECT 60.980000 61.530000 61.300000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 61.940000 61.300000 62.260000 ;
      LAYER met4 ;
        RECT 60.980000 61.940000 61.300000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 62.350000 61.300000 62.670000 ;
      LAYER met4 ;
        RECT 60.980000 62.350000 61.300000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 58.250000 61.705000 58.570000 ;
      LAYER met4 ;
        RECT 61.385000 58.250000 61.705000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 58.660000 61.705000 58.980000 ;
      LAYER met4 ;
        RECT 61.385000 58.660000 61.705000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 59.070000 61.705000 59.390000 ;
      LAYER met4 ;
        RECT 61.385000 59.070000 61.705000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 59.480000 61.705000 59.800000 ;
      LAYER met4 ;
        RECT 61.385000 59.480000 61.705000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 59.890000 61.705000 60.210000 ;
      LAYER met4 ;
        RECT 61.385000 59.890000 61.705000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 60.300000 61.705000 60.620000 ;
      LAYER met4 ;
        RECT 61.385000 60.300000 61.705000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 60.710000 61.705000 61.030000 ;
      LAYER met4 ;
        RECT 61.385000 60.710000 61.705000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 61.120000 61.705000 61.440000 ;
      LAYER met4 ;
        RECT 61.385000 61.120000 61.705000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 61.530000 61.705000 61.850000 ;
      LAYER met4 ;
        RECT 61.385000 61.530000 61.705000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 61.940000 61.705000 62.260000 ;
      LAYER met4 ;
        RECT 61.385000 61.940000 61.705000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 62.350000 61.705000 62.670000 ;
      LAYER met4 ;
        RECT 61.385000 62.350000 61.705000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 58.250000 62.110000 58.570000 ;
      LAYER met4 ;
        RECT 61.790000 58.250000 62.110000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 58.660000 62.110000 58.980000 ;
      LAYER met4 ;
        RECT 61.790000 58.660000 62.110000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 59.070000 62.110000 59.390000 ;
      LAYER met4 ;
        RECT 61.790000 59.070000 62.110000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 59.480000 62.110000 59.800000 ;
      LAYER met4 ;
        RECT 61.790000 59.480000 62.110000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 59.890000 62.110000 60.210000 ;
      LAYER met4 ;
        RECT 61.790000 59.890000 62.110000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 60.300000 62.110000 60.620000 ;
      LAYER met4 ;
        RECT 61.790000 60.300000 62.110000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 60.710000 62.110000 61.030000 ;
      LAYER met4 ;
        RECT 61.790000 60.710000 62.110000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 61.120000 62.110000 61.440000 ;
      LAYER met4 ;
        RECT 61.790000 61.120000 62.110000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 61.530000 62.110000 61.850000 ;
      LAYER met4 ;
        RECT 61.790000 61.530000 62.110000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 61.940000 62.110000 62.260000 ;
      LAYER met4 ;
        RECT 61.790000 61.940000 62.110000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 62.350000 62.110000 62.670000 ;
      LAYER met4 ;
        RECT 61.790000 62.350000 62.110000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 58.250000 62.515000 58.570000 ;
      LAYER met4 ;
        RECT 62.195000 58.250000 62.515000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 58.660000 62.515000 58.980000 ;
      LAYER met4 ;
        RECT 62.195000 58.660000 62.515000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 59.070000 62.515000 59.390000 ;
      LAYER met4 ;
        RECT 62.195000 59.070000 62.515000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 59.480000 62.515000 59.800000 ;
      LAYER met4 ;
        RECT 62.195000 59.480000 62.515000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 59.890000 62.515000 60.210000 ;
      LAYER met4 ;
        RECT 62.195000 59.890000 62.515000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 60.300000 62.515000 60.620000 ;
      LAYER met4 ;
        RECT 62.195000 60.300000 62.515000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 60.710000 62.515000 61.030000 ;
      LAYER met4 ;
        RECT 62.195000 60.710000 62.515000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 61.120000 62.515000 61.440000 ;
      LAYER met4 ;
        RECT 62.195000 61.120000 62.515000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 61.530000 62.515000 61.850000 ;
      LAYER met4 ;
        RECT 62.195000 61.530000 62.515000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 61.940000 62.515000 62.260000 ;
      LAYER met4 ;
        RECT 62.195000 61.940000 62.515000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 62.350000 62.515000 62.670000 ;
      LAYER met4 ;
        RECT 62.195000 62.350000 62.515000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 58.250000 62.920000 58.570000 ;
      LAYER met4 ;
        RECT 62.600000 58.250000 62.920000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 58.660000 62.920000 58.980000 ;
      LAYER met4 ;
        RECT 62.600000 58.660000 62.920000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 59.070000 62.920000 59.390000 ;
      LAYER met4 ;
        RECT 62.600000 59.070000 62.920000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 59.480000 62.920000 59.800000 ;
      LAYER met4 ;
        RECT 62.600000 59.480000 62.920000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 59.890000 62.920000 60.210000 ;
      LAYER met4 ;
        RECT 62.600000 59.890000 62.920000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 60.300000 62.920000 60.620000 ;
      LAYER met4 ;
        RECT 62.600000 60.300000 62.920000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 60.710000 62.920000 61.030000 ;
      LAYER met4 ;
        RECT 62.600000 60.710000 62.920000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 61.120000 62.920000 61.440000 ;
      LAYER met4 ;
        RECT 62.600000 61.120000 62.920000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 61.530000 62.920000 61.850000 ;
      LAYER met4 ;
        RECT 62.600000 61.530000 62.920000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 61.940000 62.920000 62.260000 ;
      LAYER met4 ;
        RECT 62.600000 61.940000 62.920000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 62.350000 62.920000 62.670000 ;
      LAYER met4 ;
        RECT 62.600000 62.350000 62.920000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 58.250000 63.325000 58.570000 ;
      LAYER met4 ;
        RECT 63.005000 58.250000 63.325000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 58.660000 63.325000 58.980000 ;
      LAYER met4 ;
        RECT 63.005000 58.660000 63.325000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 59.070000 63.325000 59.390000 ;
      LAYER met4 ;
        RECT 63.005000 59.070000 63.325000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 59.480000 63.325000 59.800000 ;
      LAYER met4 ;
        RECT 63.005000 59.480000 63.325000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 59.890000 63.325000 60.210000 ;
      LAYER met4 ;
        RECT 63.005000 59.890000 63.325000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 60.300000 63.325000 60.620000 ;
      LAYER met4 ;
        RECT 63.005000 60.300000 63.325000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 60.710000 63.325000 61.030000 ;
      LAYER met4 ;
        RECT 63.005000 60.710000 63.325000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 61.120000 63.325000 61.440000 ;
      LAYER met4 ;
        RECT 63.005000 61.120000 63.325000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 61.530000 63.325000 61.850000 ;
      LAYER met4 ;
        RECT 63.005000 61.530000 63.325000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 61.940000 63.325000 62.260000 ;
      LAYER met4 ;
        RECT 63.005000 61.940000 63.325000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 62.350000 63.325000 62.670000 ;
      LAYER met4 ;
        RECT 63.005000 62.350000 63.325000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 58.250000 63.730000 58.570000 ;
      LAYER met4 ;
        RECT 63.410000 58.250000 63.730000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 58.660000 63.730000 58.980000 ;
      LAYER met4 ;
        RECT 63.410000 58.660000 63.730000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 59.070000 63.730000 59.390000 ;
      LAYER met4 ;
        RECT 63.410000 59.070000 63.730000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 59.480000 63.730000 59.800000 ;
      LAYER met4 ;
        RECT 63.410000 59.480000 63.730000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 59.890000 63.730000 60.210000 ;
      LAYER met4 ;
        RECT 63.410000 59.890000 63.730000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 60.300000 63.730000 60.620000 ;
      LAYER met4 ;
        RECT 63.410000 60.300000 63.730000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 60.710000 63.730000 61.030000 ;
      LAYER met4 ;
        RECT 63.410000 60.710000 63.730000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 61.120000 63.730000 61.440000 ;
      LAYER met4 ;
        RECT 63.410000 61.120000 63.730000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 61.530000 63.730000 61.850000 ;
      LAYER met4 ;
        RECT 63.410000 61.530000 63.730000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 61.940000 63.730000 62.260000 ;
      LAYER met4 ;
        RECT 63.410000 61.940000 63.730000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 62.350000 63.730000 62.670000 ;
      LAYER met4 ;
        RECT 63.410000 62.350000 63.730000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 58.250000 64.135000 58.570000 ;
      LAYER met4 ;
        RECT 63.815000 58.250000 64.135000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 58.660000 64.135000 58.980000 ;
      LAYER met4 ;
        RECT 63.815000 58.660000 64.135000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 59.070000 64.135000 59.390000 ;
      LAYER met4 ;
        RECT 63.815000 59.070000 64.135000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 59.480000 64.135000 59.800000 ;
      LAYER met4 ;
        RECT 63.815000 59.480000 64.135000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 59.890000 64.135000 60.210000 ;
      LAYER met4 ;
        RECT 63.815000 59.890000 64.135000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 60.300000 64.135000 60.620000 ;
      LAYER met4 ;
        RECT 63.815000 60.300000 64.135000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 60.710000 64.135000 61.030000 ;
      LAYER met4 ;
        RECT 63.815000 60.710000 64.135000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 61.120000 64.135000 61.440000 ;
      LAYER met4 ;
        RECT 63.815000 61.120000 64.135000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 61.530000 64.135000 61.850000 ;
      LAYER met4 ;
        RECT 63.815000 61.530000 64.135000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 61.940000 64.135000 62.260000 ;
      LAYER met4 ;
        RECT 63.815000 61.940000 64.135000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 62.350000 64.135000 62.670000 ;
      LAYER met4 ;
        RECT 63.815000 62.350000 64.135000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 58.250000 64.540000 58.570000 ;
      LAYER met4 ;
        RECT 64.220000 58.250000 64.540000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 58.660000 64.540000 58.980000 ;
      LAYER met4 ;
        RECT 64.220000 58.660000 64.540000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 59.070000 64.540000 59.390000 ;
      LAYER met4 ;
        RECT 64.220000 59.070000 64.540000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 59.480000 64.540000 59.800000 ;
      LAYER met4 ;
        RECT 64.220000 59.480000 64.540000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 59.890000 64.540000 60.210000 ;
      LAYER met4 ;
        RECT 64.220000 59.890000 64.540000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 60.300000 64.540000 60.620000 ;
      LAYER met4 ;
        RECT 64.220000 60.300000 64.540000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 60.710000 64.540000 61.030000 ;
      LAYER met4 ;
        RECT 64.220000 60.710000 64.540000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 61.120000 64.540000 61.440000 ;
      LAYER met4 ;
        RECT 64.220000 61.120000 64.540000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 61.530000 64.540000 61.850000 ;
      LAYER met4 ;
        RECT 64.220000 61.530000 64.540000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 61.940000 64.540000 62.260000 ;
      LAYER met4 ;
        RECT 64.220000 61.940000 64.540000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 62.350000 64.540000 62.670000 ;
      LAYER met4 ;
        RECT 64.220000 62.350000 64.540000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 58.250000 64.945000 58.570000 ;
      LAYER met4 ;
        RECT 64.625000 58.250000 64.945000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 58.660000 64.945000 58.980000 ;
      LAYER met4 ;
        RECT 64.625000 58.660000 64.945000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 59.070000 64.945000 59.390000 ;
      LAYER met4 ;
        RECT 64.625000 59.070000 64.945000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 59.480000 64.945000 59.800000 ;
      LAYER met4 ;
        RECT 64.625000 59.480000 64.945000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 59.890000 64.945000 60.210000 ;
      LAYER met4 ;
        RECT 64.625000 59.890000 64.945000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 60.300000 64.945000 60.620000 ;
      LAYER met4 ;
        RECT 64.625000 60.300000 64.945000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 60.710000 64.945000 61.030000 ;
      LAYER met4 ;
        RECT 64.625000 60.710000 64.945000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 61.120000 64.945000 61.440000 ;
      LAYER met4 ;
        RECT 64.625000 61.120000 64.945000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 61.530000 64.945000 61.850000 ;
      LAYER met4 ;
        RECT 64.625000 61.530000 64.945000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 61.940000 64.945000 62.260000 ;
      LAYER met4 ;
        RECT 64.625000 61.940000 64.945000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 62.350000 64.945000 62.670000 ;
      LAYER met4 ;
        RECT 64.625000 62.350000 64.945000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 58.250000 65.350000 58.570000 ;
      LAYER met4 ;
        RECT 65.030000 58.250000 65.350000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 58.660000 65.350000 58.980000 ;
      LAYER met4 ;
        RECT 65.030000 58.660000 65.350000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 59.070000 65.350000 59.390000 ;
      LAYER met4 ;
        RECT 65.030000 59.070000 65.350000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 59.480000 65.350000 59.800000 ;
      LAYER met4 ;
        RECT 65.030000 59.480000 65.350000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 59.890000 65.350000 60.210000 ;
      LAYER met4 ;
        RECT 65.030000 59.890000 65.350000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 60.300000 65.350000 60.620000 ;
      LAYER met4 ;
        RECT 65.030000 60.300000 65.350000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 60.710000 65.350000 61.030000 ;
      LAYER met4 ;
        RECT 65.030000 60.710000 65.350000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 61.120000 65.350000 61.440000 ;
      LAYER met4 ;
        RECT 65.030000 61.120000 65.350000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 61.530000 65.350000 61.850000 ;
      LAYER met4 ;
        RECT 65.030000 61.530000 65.350000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 61.940000 65.350000 62.260000 ;
      LAYER met4 ;
        RECT 65.030000 61.940000 65.350000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 62.350000 65.350000 62.670000 ;
      LAYER met4 ;
        RECT 65.030000 62.350000 65.350000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 58.250000 65.755000 58.570000 ;
      LAYER met4 ;
        RECT 65.435000 58.250000 65.755000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 58.660000 65.755000 58.980000 ;
      LAYER met4 ;
        RECT 65.435000 58.660000 65.755000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 59.070000 65.755000 59.390000 ;
      LAYER met4 ;
        RECT 65.435000 59.070000 65.755000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 59.480000 65.755000 59.800000 ;
      LAYER met4 ;
        RECT 65.435000 59.480000 65.755000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 59.890000 65.755000 60.210000 ;
      LAYER met4 ;
        RECT 65.435000 59.890000 65.755000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 60.300000 65.755000 60.620000 ;
      LAYER met4 ;
        RECT 65.435000 60.300000 65.755000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 60.710000 65.755000 61.030000 ;
      LAYER met4 ;
        RECT 65.435000 60.710000 65.755000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 61.120000 65.755000 61.440000 ;
      LAYER met4 ;
        RECT 65.435000 61.120000 65.755000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 61.530000 65.755000 61.850000 ;
      LAYER met4 ;
        RECT 65.435000 61.530000 65.755000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 61.940000 65.755000 62.260000 ;
      LAYER met4 ;
        RECT 65.435000 61.940000 65.755000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 62.350000 65.755000 62.670000 ;
      LAYER met4 ;
        RECT 65.435000 62.350000 65.755000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 58.250000 66.160000 58.570000 ;
      LAYER met4 ;
        RECT 65.840000 58.250000 66.160000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 58.660000 66.160000 58.980000 ;
      LAYER met4 ;
        RECT 65.840000 58.660000 66.160000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 59.070000 66.160000 59.390000 ;
      LAYER met4 ;
        RECT 65.840000 59.070000 66.160000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 59.480000 66.160000 59.800000 ;
      LAYER met4 ;
        RECT 65.840000 59.480000 66.160000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 59.890000 66.160000 60.210000 ;
      LAYER met4 ;
        RECT 65.840000 59.890000 66.160000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 60.300000 66.160000 60.620000 ;
      LAYER met4 ;
        RECT 65.840000 60.300000 66.160000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 60.710000 66.160000 61.030000 ;
      LAYER met4 ;
        RECT 65.840000 60.710000 66.160000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 61.120000 66.160000 61.440000 ;
      LAYER met4 ;
        RECT 65.840000 61.120000 66.160000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 61.530000 66.160000 61.850000 ;
      LAYER met4 ;
        RECT 65.840000 61.530000 66.160000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 61.940000 66.160000 62.260000 ;
      LAYER met4 ;
        RECT 65.840000 61.940000 66.160000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 62.350000 66.160000 62.670000 ;
      LAYER met4 ;
        RECT 65.840000 62.350000 66.160000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 58.250000 66.565000 58.570000 ;
      LAYER met4 ;
        RECT 66.245000 58.250000 66.565000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 58.660000 66.565000 58.980000 ;
      LAYER met4 ;
        RECT 66.245000 58.660000 66.565000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 59.070000 66.565000 59.390000 ;
      LAYER met4 ;
        RECT 66.245000 59.070000 66.565000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 59.480000 66.565000 59.800000 ;
      LAYER met4 ;
        RECT 66.245000 59.480000 66.565000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 59.890000 66.565000 60.210000 ;
      LAYER met4 ;
        RECT 66.245000 59.890000 66.565000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 60.300000 66.565000 60.620000 ;
      LAYER met4 ;
        RECT 66.245000 60.300000 66.565000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 60.710000 66.565000 61.030000 ;
      LAYER met4 ;
        RECT 66.245000 60.710000 66.565000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 61.120000 66.565000 61.440000 ;
      LAYER met4 ;
        RECT 66.245000 61.120000 66.565000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 61.530000 66.565000 61.850000 ;
      LAYER met4 ;
        RECT 66.245000 61.530000 66.565000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 61.940000 66.565000 62.260000 ;
      LAYER met4 ;
        RECT 66.245000 61.940000 66.565000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 62.350000 66.565000 62.670000 ;
      LAYER met4 ;
        RECT 66.245000 62.350000 66.565000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 58.250000 66.970000 58.570000 ;
      LAYER met4 ;
        RECT 66.650000 58.250000 66.970000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 58.660000 66.970000 58.980000 ;
      LAYER met4 ;
        RECT 66.650000 58.660000 66.970000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 59.070000 66.970000 59.390000 ;
      LAYER met4 ;
        RECT 66.650000 59.070000 66.970000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 59.480000 66.970000 59.800000 ;
      LAYER met4 ;
        RECT 66.650000 59.480000 66.970000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 59.890000 66.970000 60.210000 ;
      LAYER met4 ;
        RECT 66.650000 59.890000 66.970000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 60.300000 66.970000 60.620000 ;
      LAYER met4 ;
        RECT 66.650000 60.300000 66.970000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 60.710000 66.970000 61.030000 ;
      LAYER met4 ;
        RECT 66.650000 60.710000 66.970000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 61.120000 66.970000 61.440000 ;
      LAYER met4 ;
        RECT 66.650000 61.120000 66.970000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 61.530000 66.970000 61.850000 ;
      LAYER met4 ;
        RECT 66.650000 61.530000 66.970000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 61.940000 66.970000 62.260000 ;
      LAYER met4 ;
        RECT 66.650000 61.940000 66.970000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 62.350000 66.970000 62.670000 ;
      LAYER met4 ;
        RECT 66.650000 62.350000 66.970000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 58.250000 67.375000 58.570000 ;
      LAYER met4 ;
        RECT 67.055000 58.250000 67.375000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 58.660000 67.375000 58.980000 ;
      LAYER met4 ;
        RECT 67.055000 58.660000 67.375000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 59.070000 67.375000 59.390000 ;
      LAYER met4 ;
        RECT 67.055000 59.070000 67.375000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 59.480000 67.375000 59.800000 ;
      LAYER met4 ;
        RECT 67.055000 59.480000 67.375000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 59.890000 67.375000 60.210000 ;
      LAYER met4 ;
        RECT 67.055000 59.890000 67.375000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 60.300000 67.375000 60.620000 ;
      LAYER met4 ;
        RECT 67.055000 60.300000 67.375000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 60.710000 67.375000 61.030000 ;
      LAYER met4 ;
        RECT 67.055000 60.710000 67.375000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 61.120000 67.375000 61.440000 ;
      LAYER met4 ;
        RECT 67.055000 61.120000 67.375000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 61.530000 67.375000 61.850000 ;
      LAYER met4 ;
        RECT 67.055000 61.530000 67.375000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 61.940000 67.375000 62.260000 ;
      LAYER met4 ;
        RECT 67.055000 61.940000 67.375000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 62.350000 67.375000 62.670000 ;
      LAYER met4 ;
        RECT 67.055000 62.350000 67.375000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 58.250000 67.780000 58.570000 ;
      LAYER met4 ;
        RECT 67.460000 58.250000 67.780000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 58.660000 67.780000 58.980000 ;
      LAYER met4 ;
        RECT 67.460000 58.660000 67.780000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 59.070000 67.780000 59.390000 ;
      LAYER met4 ;
        RECT 67.460000 59.070000 67.780000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 59.480000 67.780000 59.800000 ;
      LAYER met4 ;
        RECT 67.460000 59.480000 67.780000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 59.890000 67.780000 60.210000 ;
      LAYER met4 ;
        RECT 67.460000 59.890000 67.780000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 60.300000 67.780000 60.620000 ;
      LAYER met4 ;
        RECT 67.460000 60.300000 67.780000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 60.710000 67.780000 61.030000 ;
      LAYER met4 ;
        RECT 67.460000 60.710000 67.780000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 61.120000 67.780000 61.440000 ;
      LAYER met4 ;
        RECT 67.460000 61.120000 67.780000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 61.530000 67.780000 61.850000 ;
      LAYER met4 ;
        RECT 67.460000 61.530000 67.780000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 61.940000 67.780000 62.260000 ;
      LAYER met4 ;
        RECT 67.460000 61.940000 67.780000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 62.350000 67.780000 62.670000 ;
      LAYER met4 ;
        RECT 67.460000 62.350000 67.780000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 58.250000 68.185000 58.570000 ;
      LAYER met4 ;
        RECT 67.865000 58.250000 68.185000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 58.660000 68.185000 58.980000 ;
      LAYER met4 ;
        RECT 67.865000 58.660000 68.185000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 59.070000 68.185000 59.390000 ;
      LAYER met4 ;
        RECT 67.865000 59.070000 68.185000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 59.480000 68.185000 59.800000 ;
      LAYER met4 ;
        RECT 67.865000 59.480000 68.185000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 59.890000 68.185000 60.210000 ;
      LAYER met4 ;
        RECT 67.865000 59.890000 68.185000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 60.300000 68.185000 60.620000 ;
      LAYER met4 ;
        RECT 67.865000 60.300000 68.185000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 60.710000 68.185000 61.030000 ;
      LAYER met4 ;
        RECT 67.865000 60.710000 68.185000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 61.120000 68.185000 61.440000 ;
      LAYER met4 ;
        RECT 67.865000 61.120000 68.185000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 61.530000 68.185000 61.850000 ;
      LAYER met4 ;
        RECT 67.865000 61.530000 68.185000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 61.940000 68.185000 62.260000 ;
      LAYER met4 ;
        RECT 67.865000 61.940000 68.185000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 62.350000 68.185000 62.670000 ;
      LAYER met4 ;
        RECT 67.865000 62.350000 68.185000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 58.250000 68.590000 58.570000 ;
      LAYER met4 ;
        RECT 68.270000 58.250000 68.590000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 58.660000 68.590000 58.980000 ;
      LAYER met4 ;
        RECT 68.270000 58.660000 68.590000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 59.070000 68.590000 59.390000 ;
      LAYER met4 ;
        RECT 68.270000 59.070000 68.590000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 59.480000 68.590000 59.800000 ;
      LAYER met4 ;
        RECT 68.270000 59.480000 68.590000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 59.890000 68.590000 60.210000 ;
      LAYER met4 ;
        RECT 68.270000 59.890000 68.590000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 60.300000 68.590000 60.620000 ;
      LAYER met4 ;
        RECT 68.270000 60.300000 68.590000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 60.710000 68.590000 61.030000 ;
      LAYER met4 ;
        RECT 68.270000 60.710000 68.590000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 61.120000 68.590000 61.440000 ;
      LAYER met4 ;
        RECT 68.270000 61.120000 68.590000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 61.530000 68.590000 61.850000 ;
      LAYER met4 ;
        RECT 68.270000 61.530000 68.590000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 61.940000 68.590000 62.260000 ;
      LAYER met4 ;
        RECT 68.270000 61.940000 68.590000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 62.350000 68.590000 62.670000 ;
      LAYER met4 ;
        RECT 68.270000 62.350000 68.590000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 58.250000 68.995000 58.570000 ;
      LAYER met4 ;
        RECT 68.675000 58.250000 68.995000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 58.660000 68.995000 58.980000 ;
      LAYER met4 ;
        RECT 68.675000 58.660000 68.995000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 59.070000 68.995000 59.390000 ;
      LAYER met4 ;
        RECT 68.675000 59.070000 68.995000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 59.480000 68.995000 59.800000 ;
      LAYER met4 ;
        RECT 68.675000 59.480000 68.995000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 59.890000 68.995000 60.210000 ;
      LAYER met4 ;
        RECT 68.675000 59.890000 68.995000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 60.300000 68.995000 60.620000 ;
      LAYER met4 ;
        RECT 68.675000 60.300000 68.995000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 60.710000 68.995000 61.030000 ;
      LAYER met4 ;
        RECT 68.675000 60.710000 68.995000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 61.120000 68.995000 61.440000 ;
      LAYER met4 ;
        RECT 68.675000 61.120000 68.995000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 61.530000 68.995000 61.850000 ;
      LAYER met4 ;
        RECT 68.675000 61.530000 68.995000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 61.940000 68.995000 62.260000 ;
      LAYER met4 ;
        RECT 68.675000 61.940000 68.995000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 62.350000 68.995000 62.670000 ;
      LAYER met4 ;
        RECT 68.675000 62.350000 68.995000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 58.250000 69.400000 58.570000 ;
      LAYER met4 ;
        RECT 69.080000 58.250000 69.400000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 58.660000 69.400000 58.980000 ;
      LAYER met4 ;
        RECT 69.080000 58.660000 69.400000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 59.070000 69.400000 59.390000 ;
      LAYER met4 ;
        RECT 69.080000 59.070000 69.400000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 59.480000 69.400000 59.800000 ;
      LAYER met4 ;
        RECT 69.080000 59.480000 69.400000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 59.890000 69.400000 60.210000 ;
      LAYER met4 ;
        RECT 69.080000 59.890000 69.400000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 60.300000 69.400000 60.620000 ;
      LAYER met4 ;
        RECT 69.080000 60.300000 69.400000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 60.710000 69.400000 61.030000 ;
      LAYER met4 ;
        RECT 69.080000 60.710000 69.400000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 61.120000 69.400000 61.440000 ;
      LAYER met4 ;
        RECT 69.080000 61.120000 69.400000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 61.530000 69.400000 61.850000 ;
      LAYER met4 ;
        RECT 69.080000 61.530000 69.400000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 61.940000 69.400000 62.260000 ;
      LAYER met4 ;
        RECT 69.080000 61.940000 69.400000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 62.350000 69.400000 62.670000 ;
      LAYER met4 ;
        RECT 69.080000 62.350000 69.400000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 58.250000 69.805000 58.570000 ;
      LAYER met4 ;
        RECT 69.485000 58.250000 69.805000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 58.660000 69.805000 58.980000 ;
      LAYER met4 ;
        RECT 69.485000 58.660000 69.805000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 59.070000 69.805000 59.390000 ;
      LAYER met4 ;
        RECT 69.485000 59.070000 69.805000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 59.480000 69.805000 59.800000 ;
      LAYER met4 ;
        RECT 69.485000 59.480000 69.805000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 59.890000 69.805000 60.210000 ;
      LAYER met4 ;
        RECT 69.485000 59.890000 69.805000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 60.300000 69.805000 60.620000 ;
      LAYER met4 ;
        RECT 69.485000 60.300000 69.805000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 60.710000 69.805000 61.030000 ;
      LAYER met4 ;
        RECT 69.485000 60.710000 69.805000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 61.120000 69.805000 61.440000 ;
      LAYER met4 ;
        RECT 69.485000 61.120000 69.805000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 61.530000 69.805000 61.850000 ;
      LAYER met4 ;
        RECT 69.485000 61.530000 69.805000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 61.940000 69.805000 62.260000 ;
      LAYER met4 ;
        RECT 69.485000 61.940000 69.805000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 62.350000 69.805000 62.670000 ;
      LAYER met4 ;
        RECT 69.485000 62.350000 69.805000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 58.250000 70.210000 58.570000 ;
      LAYER met4 ;
        RECT 69.890000 58.250000 70.210000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 58.660000 70.210000 58.980000 ;
      LAYER met4 ;
        RECT 69.890000 58.660000 70.210000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 59.070000 70.210000 59.390000 ;
      LAYER met4 ;
        RECT 69.890000 59.070000 70.210000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 59.480000 70.210000 59.800000 ;
      LAYER met4 ;
        RECT 69.890000 59.480000 70.210000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 59.890000 70.210000 60.210000 ;
      LAYER met4 ;
        RECT 69.890000 59.890000 70.210000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 60.300000 70.210000 60.620000 ;
      LAYER met4 ;
        RECT 69.890000 60.300000 70.210000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 60.710000 70.210000 61.030000 ;
      LAYER met4 ;
        RECT 69.890000 60.710000 70.210000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 61.120000 70.210000 61.440000 ;
      LAYER met4 ;
        RECT 69.890000 61.120000 70.210000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 61.530000 70.210000 61.850000 ;
      LAYER met4 ;
        RECT 69.890000 61.530000 70.210000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 61.940000 70.210000 62.260000 ;
      LAYER met4 ;
        RECT 69.890000 61.940000 70.210000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 62.350000 70.210000 62.670000 ;
      LAYER met4 ;
        RECT 69.890000 62.350000 70.210000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 58.250000 7.355000 58.570000 ;
      LAYER met4 ;
        RECT 7.035000 58.250000 7.355000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 58.660000 7.355000 58.980000 ;
      LAYER met4 ;
        RECT 7.035000 58.660000 7.355000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 59.070000 7.355000 59.390000 ;
      LAYER met4 ;
        RECT 7.035000 59.070000 7.355000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 59.480000 7.355000 59.800000 ;
      LAYER met4 ;
        RECT 7.035000 59.480000 7.355000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 59.890000 7.355000 60.210000 ;
      LAYER met4 ;
        RECT 7.035000 59.890000 7.355000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 60.300000 7.355000 60.620000 ;
      LAYER met4 ;
        RECT 7.035000 60.300000 7.355000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 60.710000 7.355000 61.030000 ;
      LAYER met4 ;
        RECT 7.035000 60.710000 7.355000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 61.120000 7.355000 61.440000 ;
      LAYER met4 ;
        RECT 7.035000 61.120000 7.355000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 61.530000 7.355000 61.850000 ;
      LAYER met4 ;
        RECT 7.035000 61.530000 7.355000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 61.940000 7.355000 62.260000 ;
      LAYER met4 ;
        RECT 7.035000 61.940000 7.355000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 62.350000 7.355000 62.670000 ;
      LAYER met4 ;
        RECT 7.035000 62.350000 7.355000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 58.250000 7.760000 58.570000 ;
      LAYER met4 ;
        RECT 7.440000 58.250000 7.760000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 58.660000 7.760000 58.980000 ;
      LAYER met4 ;
        RECT 7.440000 58.660000 7.760000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 59.070000 7.760000 59.390000 ;
      LAYER met4 ;
        RECT 7.440000 59.070000 7.760000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 59.480000 7.760000 59.800000 ;
      LAYER met4 ;
        RECT 7.440000 59.480000 7.760000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 59.890000 7.760000 60.210000 ;
      LAYER met4 ;
        RECT 7.440000 59.890000 7.760000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 60.300000 7.760000 60.620000 ;
      LAYER met4 ;
        RECT 7.440000 60.300000 7.760000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 60.710000 7.760000 61.030000 ;
      LAYER met4 ;
        RECT 7.440000 60.710000 7.760000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 61.120000 7.760000 61.440000 ;
      LAYER met4 ;
        RECT 7.440000 61.120000 7.760000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 61.530000 7.760000 61.850000 ;
      LAYER met4 ;
        RECT 7.440000 61.530000 7.760000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 61.940000 7.760000 62.260000 ;
      LAYER met4 ;
        RECT 7.440000 61.940000 7.760000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 62.350000 7.760000 62.670000 ;
      LAYER met4 ;
        RECT 7.440000 62.350000 7.760000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 58.250000 8.165000 58.570000 ;
      LAYER met4 ;
        RECT 7.845000 58.250000 8.165000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 58.660000 8.165000 58.980000 ;
      LAYER met4 ;
        RECT 7.845000 58.660000 8.165000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 59.070000 8.165000 59.390000 ;
      LAYER met4 ;
        RECT 7.845000 59.070000 8.165000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 59.480000 8.165000 59.800000 ;
      LAYER met4 ;
        RECT 7.845000 59.480000 8.165000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 59.890000 8.165000 60.210000 ;
      LAYER met4 ;
        RECT 7.845000 59.890000 8.165000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 60.300000 8.165000 60.620000 ;
      LAYER met4 ;
        RECT 7.845000 60.300000 8.165000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 60.710000 8.165000 61.030000 ;
      LAYER met4 ;
        RECT 7.845000 60.710000 8.165000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 61.120000 8.165000 61.440000 ;
      LAYER met4 ;
        RECT 7.845000 61.120000 8.165000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 61.530000 8.165000 61.850000 ;
      LAYER met4 ;
        RECT 7.845000 61.530000 8.165000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 61.940000 8.165000 62.260000 ;
      LAYER met4 ;
        RECT 7.845000 61.940000 8.165000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 62.350000 8.165000 62.670000 ;
      LAYER met4 ;
        RECT 7.845000 62.350000 8.165000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 58.250000 70.615000 58.570000 ;
      LAYER met4 ;
        RECT 70.295000 58.250000 70.615000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 58.660000 70.615000 58.980000 ;
      LAYER met4 ;
        RECT 70.295000 58.660000 70.615000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 59.070000 70.615000 59.390000 ;
      LAYER met4 ;
        RECT 70.295000 59.070000 70.615000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 59.480000 70.615000 59.800000 ;
      LAYER met4 ;
        RECT 70.295000 59.480000 70.615000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 59.890000 70.615000 60.210000 ;
      LAYER met4 ;
        RECT 70.295000 59.890000 70.615000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 60.300000 70.615000 60.620000 ;
      LAYER met4 ;
        RECT 70.295000 60.300000 70.615000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 60.710000 70.615000 61.030000 ;
      LAYER met4 ;
        RECT 70.295000 60.710000 70.615000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 61.120000 70.615000 61.440000 ;
      LAYER met4 ;
        RECT 70.295000 61.120000 70.615000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 61.530000 70.615000 61.850000 ;
      LAYER met4 ;
        RECT 70.295000 61.530000 70.615000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 61.940000 70.615000 62.260000 ;
      LAYER met4 ;
        RECT 70.295000 61.940000 70.615000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 62.350000 70.615000 62.670000 ;
      LAYER met4 ;
        RECT 70.295000 62.350000 70.615000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 58.250000 71.020000 58.570000 ;
      LAYER met4 ;
        RECT 70.700000 58.250000 71.020000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 58.660000 71.020000 58.980000 ;
      LAYER met4 ;
        RECT 70.700000 58.660000 71.020000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 59.070000 71.020000 59.390000 ;
      LAYER met4 ;
        RECT 70.700000 59.070000 71.020000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 59.480000 71.020000 59.800000 ;
      LAYER met4 ;
        RECT 70.700000 59.480000 71.020000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 59.890000 71.020000 60.210000 ;
      LAYER met4 ;
        RECT 70.700000 59.890000 71.020000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 60.300000 71.020000 60.620000 ;
      LAYER met4 ;
        RECT 70.700000 60.300000 71.020000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 60.710000 71.020000 61.030000 ;
      LAYER met4 ;
        RECT 70.700000 60.710000 71.020000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 61.120000 71.020000 61.440000 ;
      LAYER met4 ;
        RECT 70.700000 61.120000 71.020000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 61.530000 71.020000 61.850000 ;
      LAYER met4 ;
        RECT 70.700000 61.530000 71.020000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 61.940000 71.020000 62.260000 ;
      LAYER met4 ;
        RECT 70.700000 61.940000 71.020000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 62.350000 71.020000 62.670000 ;
      LAYER met4 ;
        RECT 70.700000 62.350000 71.020000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 58.250000 71.425000 58.570000 ;
      LAYER met4 ;
        RECT 71.105000 58.250000 71.425000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 58.660000 71.425000 58.980000 ;
      LAYER met4 ;
        RECT 71.105000 58.660000 71.425000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 59.070000 71.425000 59.390000 ;
      LAYER met4 ;
        RECT 71.105000 59.070000 71.425000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 59.480000 71.425000 59.800000 ;
      LAYER met4 ;
        RECT 71.105000 59.480000 71.425000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 59.890000 71.425000 60.210000 ;
      LAYER met4 ;
        RECT 71.105000 59.890000 71.425000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 60.300000 71.425000 60.620000 ;
      LAYER met4 ;
        RECT 71.105000 60.300000 71.425000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 60.710000 71.425000 61.030000 ;
      LAYER met4 ;
        RECT 71.105000 60.710000 71.425000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 61.120000 71.425000 61.440000 ;
      LAYER met4 ;
        RECT 71.105000 61.120000 71.425000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 61.530000 71.425000 61.850000 ;
      LAYER met4 ;
        RECT 71.105000 61.530000 71.425000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 61.940000 71.425000 62.260000 ;
      LAYER met4 ;
        RECT 71.105000 61.940000 71.425000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 62.350000 71.425000 62.670000 ;
      LAYER met4 ;
        RECT 71.105000 62.350000 71.425000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 58.250000 71.830000 58.570000 ;
      LAYER met4 ;
        RECT 71.510000 58.250000 71.830000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 58.660000 71.830000 58.980000 ;
      LAYER met4 ;
        RECT 71.510000 58.660000 71.830000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 59.070000 71.830000 59.390000 ;
      LAYER met4 ;
        RECT 71.510000 59.070000 71.830000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 59.480000 71.830000 59.800000 ;
      LAYER met4 ;
        RECT 71.510000 59.480000 71.830000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 59.890000 71.830000 60.210000 ;
      LAYER met4 ;
        RECT 71.510000 59.890000 71.830000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 60.300000 71.830000 60.620000 ;
      LAYER met4 ;
        RECT 71.510000 60.300000 71.830000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 60.710000 71.830000 61.030000 ;
      LAYER met4 ;
        RECT 71.510000 60.710000 71.830000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 61.120000 71.830000 61.440000 ;
      LAYER met4 ;
        RECT 71.510000 61.120000 71.830000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 61.530000 71.830000 61.850000 ;
      LAYER met4 ;
        RECT 71.510000 61.530000 71.830000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 61.940000 71.830000 62.260000 ;
      LAYER met4 ;
        RECT 71.510000 61.940000 71.830000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 62.350000 71.830000 62.670000 ;
      LAYER met4 ;
        RECT 71.510000 62.350000 71.830000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 58.250000 72.235000 58.570000 ;
      LAYER met4 ;
        RECT 71.915000 58.250000 72.235000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 58.660000 72.235000 58.980000 ;
      LAYER met4 ;
        RECT 71.915000 58.660000 72.235000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 59.070000 72.235000 59.390000 ;
      LAYER met4 ;
        RECT 71.915000 59.070000 72.235000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 59.480000 72.235000 59.800000 ;
      LAYER met4 ;
        RECT 71.915000 59.480000 72.235000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 59.890000 72.235000 60.210000 ;
      LAYER met4 ;
        RECT 71.915000 59.890000 72.235000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 60.300000 72.235000 60.620000 ;
      LAYER met4 ;
        RECT 71.915000 60.300000 72.235000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 60.710000 72.235000 61.030000 ;
      LAYER met4 ;
        RECT 71.915000 60.710000 72.235000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 61.120000 72.235000 61.440000 ;
      LAYER met4 ;
        RECT 71.915000 61.120000 72.235000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 61.530000 72.235000 61.850000 ;
      LAYER met4 ;
        RECT 71.915000 61.530000 72.235000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 61.940000 72.235000 62.260000 ;
      LAYER met4 ;
        RECT 71.915000 61.940000 72.235000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 62.350000 72.235000 62.670000 ;
      LAYER met4 ;
        RECT 71.915000 62.350000 72.235000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 58.250000 72.640000 58.570000 ;
      LAYER met4 ;
        RECT 72.320000 58.250000 72.640000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 58.660000 72.640000 58.980000 ;
      LAYER met4 ;
        RECT 72.320000 58.660000 72.640000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 59.070000 72.640000 59.390000 ;
      LAYER met4 ;
        RECT 72.320000 59.070000 72.640000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 59.480000 72.640000 59.800000 ;
      LAYER met4 ;
        RECT 72.320000 59.480000 72.640000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 59.890000 72.640000 60.210000 ;
      LAYER met4 ;
        RECT 72.320000 59.890000 72.640000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 60.300000 72.640000 60.620000 ;
      LAYER met4 ;
        RECT 72.320000 60.300000 72.640000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 60.710000 72.640000 61.030000 ;
      LAYER met4 ;
        RECT 72.320000 60.710000 72.640000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 61.120000 72.640000 61.440000 ;
      LAYER met4 ;
        RECT 72.320000 61.120000 72.640000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 61.530000 72.640000 61.850000 ;
      LAYER met4 ;
        RECT 72.320000 61.530000 72.640000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 61.940000 72.640000 62.260000 ;
      LAYER met4 ;
        RECT 72.320000 61.940000 72.640000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 62.350000 72.640000 62.670000 ;
      LAYER met4 ;
        RECT 72.320000 62.350000 72.640000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 58.250000 73.045000 58.570000 ;
      LAYER met4 ;
        RECT 72.725000 58.250000 73.045000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 58.660000 73.045000 58.980000 ;
      LAYER met4 ;
        RECT 72.725000 58.660000 73.045000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 59.070000 73.045000 59.390000 ;
      LAYER met4 ;
        RECT 72.725000 59.070000 73.045000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 59.480000 73.045000 59.800000 ;
      LAYER met4 ;
        RECT 72.725000 59.480000 73.045000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 59.890000 73.045000 60.210000 ;
      LAYER met4 ;
        RECT 72.725000 59.890000 73.045000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 60.300000 73.045000 60.620000 ;
      LAYER met4 ;
        RECT 72.725000 60.300000 73.045000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 60.710000 73.045000 61.030000 ;
      LAYER met4 ;
        RECT 72.725000 60.710000 73.045000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 61.120000 73.045000 61.440000 ;
      LAYER met4 ;
        RECT 72.725000 61.120000 73.045000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 61.530000 73.045000 61.850000 ;
      LAYER met4 ;
        RECT 72.725000 61.530000 73.045000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 61.940000 73.045000 62.260000 ;
      LAYER met4 ;
        RECT 72.725000 61.940000 73.045000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 62.350000 73.045000 62.670000 ;
      LAYER met4 ;
        RECT 72.725000 62.350000 73.045000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 58.250000 73.450000 58.570000 ;
      LAYER met4 ;
        RECT 73.130000 58.250000 73.450000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 58.660000 73.450000 58.980000 ;
      LAYER met4 ;
        RECT 73.130000 58.660000 73.450000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 59.070000 73.450000 59.390000 ;
      LAYER met4 ;
        RECT 73.130000 59.070000 73.450000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 59.480000 73.450000 59.800000 ;
      LAYER met4 ;
        RECT 73.130000 59.480000 73.450000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 59.890000 73.450000 60.210000 ;
      LAYER met4 ;
        RECT 73.130000 59.890000 73.450000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 60.300000 73.450000 60.620000 ;
      LAYER met4 ;
        RECT 73.130000 60.300000 73.450000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 60.710000 73.450000 61.030000 ;
      LAYER met4 ;
        RECT 73.130000 60.710000 73.450000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 61.120000 73.450000 61.440000 ;
      LAYER met4 ;
        RECT 73.130000 61.120000 73.450000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 61.530000 73.450000 61.850000 ;
      LAYER met4 ;
        RECT 73.130000 61.530000 73.450000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 61.940000 73.450000 62.260000 ;
      LAYER met4 ;
        RECT 73.130000 61.940000 73.450000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 62.350000 73.450000 62.670000 ;
      LAYER met4 ;
        RECT 73.130000 62.350000 73.450000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 58.250000 73.855000 58.570000 ;
      LAYER met4 ;
        RECT 73.535000 58.250000 73.855000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 58.660000 73.855000 58.980000 ;
      LAYER met4 ;
        RECT 73.535000 58.660000 73.855000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 59.070000 73.855000 59.390000 ;
      LAYER met4 ;
        RECT 73.535000 59.070000 73.855000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 59.480000 73.855000 59.800000 ;
      LAYER met4 ;
        RECT 73.535000 59.480000 73.855000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 59.890000 73.855000 60.210000 ;
      LAYER met4 ;
        RECT 73.535000 59.890000 73.855000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 60.300000 73.855000 60.620000 ;
      LAYER met4 ;
        RECT 73.535000 60.300000 73.855000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 60.710000 73.855000 61.030000 ;
      LAYER met4 ;
        RECT 73.535000 60.710000 73.855000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 61.120000 73.855000 61.440000 ;
      LAYER met4 ;
        RECT 73.535000 61.120000 73.855000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 61.530000 73.855000 61.850000 ;
      LAYER met4 ;
        RECT 73.535000 61.530000 73.855000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 61.940000 73.855000 62.260000 ;
      LAYER met4 ;
        RECT 73.535000 61.940000 73.855000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 62.350000 73.855000 62.670000 ;
      LAYER met4 ;
        RECT 73.535000 62.350000 73.855000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 58.250000 74.260000 58.570000 ;
      LAYER met4 ;
        RECT 73.940000 58.250000 74.260000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 58.660000 74.260000 58.980000 ;
      LAYER met4 ;
        RECT 73.940000 58.660000 74.260000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 59.070000 74.260000 59.390000 ;
      LAYER met4 ;
        RECT 73.940000 59.070000 74.260000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 59.480000 74.260000 59.800000 ;
      LAYER met4 ;
        RECT 73.940000 59.480000 74.260000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 59.890000 74.260000 60.210000 ;
      LAYER met4 ;
        RECT 73.940000 59.890000 74.260000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 60.300000 74.260000 60.620000 ;
      LAYER met4 ;
        RECT 73.940000 60.300000 74.260000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 60.710000 74.260000 61.030000 ;
      LAYER met4 ;
        RECT 73.940000 60.710000 74.260000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 61.120000 74.260000 61.440000 ;
      LAYER met4 ;
        RECT 73.940000 61.120000 74.260000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 61.530000 74.260000 61.850000 ;
      LAYER met4 ;
        RECT 73.940000 61.530000 74.260000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 61.940000 74.260000 62.260000 ;
      LAYER met4 ;
        RECT 73.940000 61.940000 74.260000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 62.350000 74.260000 62.670000 ;
      LAYER met4 ;
        RECT 73.940000 62.350000 74.260000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 58.250000 8.570000 58.570000 ;
      LAYER met4 ;
        RECT 8.250000 58.250000 8.570000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 58.660000 8.570000 58.980000 ;
      LAYER met4 ;
        RECT 8.250000 58.660000 8.570000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 59.070000 8.570000 59.390000 ;
      LAYER met4 ;
        RECT 8.250000 59.070000 8.570000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 59.480000 8.570000 59.800000 ;
      LAYER met4 ;
        RECT 8.250000 59.480000 8.570000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 59.890000 8.570000 60.210000 ;
      LAYER met4 ;
        RECT 8.250000 59.890000 8.570000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 60.300000 8.570000 60.620000 ;
      LAYER met4 ;
        RECT 8.250000 60.300000 8.570000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 60.710000 8.570000 61.030000 ;
      LAYER met4 ;
        RECT 8.250000 60.710000 8.570000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 61.120000 8.570000 61.440000 ;
      LAYER met4 ;
        RECT 8.250000 61.120000 8.570000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 61.530000 8.570000 61.850000 ;
      LAYER met4 ;
        RECT 8.250000 61.530000 8.570000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 61.940000 8.570000 62.260000 ;
      LAYER met4 ;
        RECT 8.250000 61.940000 8.570000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 62.350000 8.570000 62.670000 ;
      LAYER met4 ;
        RECT 8.250000 62.350000 8.570000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 58.250000 8.975000 58.570000 ;
      LAYER met4 ;
        RECT 8.655000 58.250000 8.975000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 58.660000 8.975000 58.980000 ;
      LAYER met4 ;
        RECT 8.655000 58.660000 8.975000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 59.070000 8.975000 59.390000 ;
      LAYER met4 ;
        RECT 8.655000 59.070000 8.975000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 59.480000 8.975000 59.800000 ;
      LAYER met4 ;
        RECT 8.655000 59.480000 8.975000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 59.890000 8.975000 60.210000 ;
      LAYER met4 ;
        RECT 8.655000 59.890000 8.975000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 60.300000 8.975000 60.620000 ;
      LAYER met4 ;
        RECT 8.655000 60.300000 8.975000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 60.710000 8.975000 61.030000 ;
      LAYER met4 ;
        RECT 8.655000 60.710000 8.975000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 61.120000 8.975000 61.440000 ;
      LAYER met4 ;
        RECT 8.655000 61.120000 8.975000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 61.530000 8.975000 61.850000 ;
      LAYER met4 ;
        RECT 8.655000 61.530000 8.975000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 61.940000 8.975000 62.260000 ;
      LAYER met4 ;
        RECT 8.655000 61.940000 8.975000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 62.350000 8.975000 62.670000 ;
      LAYER met4 ;
        RECT 8.655000 62.350000 8.975000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 58.250000 9.380000 58.570000 ;
      LAYER met4 ;
        RECT 9.060000 58.250000 9.380000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 58.660000 9.380000 58.980000 ;
      LAYER met4 ;
        RECT 9.060000 58.660000 9.380000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 59.070000 9.380000 59.390000 ;
      LAYER met4 ;
        RECT 9.060000 59.070000 9.380000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 59.480000 9.380000 59.800000 ;
      LAYER met4 ;
        RECT 9.060000 59.480000 9.380000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 59.890000 9.380000 60.210000 ;
      LAYER met4 ;
        RECT 9.060000 59.890000 9.380000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 60.300000 9.380000 60.620000 ;
      LAYER met4 ;
        RECT 9.060000 60.300000 9.380000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 60.710000 9.380000 61.030000 ;
      LAYER met4 ;
        RECT 9.060000 60.710000 9.380000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 61.120000 9.380000 61.440000 ;
      LAYER met4 ;
        RECT 9.060000 61.120000 9.380000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 61.530000 9.380000 61.850000 ;
      LAYER met4 ;
        RECT 9.060000 61.530000 9.380000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 61.940000 9.380000 62.260000 ;
      LAYER met4 ;
        RECT 9.060000 61.940000 9.380000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 62.350000 9.380000 62.670000 ;
      LAYER met4 ;
        RECT 9.060000 62.350000 9.380000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 58.250000 9.785000 58.570000 ;
      LAYER met4 ;
        RECT 9.465000 58.250000 9.785000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 58.660000 9.785000 58.980000 ;
      LAYER met4 ;
        RECT 9.465000 58.660000 9.785000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 59.070000 9.785000 59.390000 ;
      LAYER met4 ;
        RECT 9.465000 59.070000 9.785000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 59.480000 9.785000 59.800000 ;
      LAYER met4 ;
        RECT 9.465000 59.480000 9.785000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 59.890000 9.785000 60.210000 ;
      LAYER met4 ;
        RECT 9.465000 59.890000 9.785000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 60.300000 9.785000 60.620000 ;
      LAYER met4 ;
        RECT 9.465000 60.300000 9.785000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 60.710000 9.785000 61.030000 ;
      LAYER met4 ;
        RECT 9.465000 60.710000 9.785000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 61.120000 9.785000 61.440000 ;
      LAYER met4 ;
        RECT 9.465000 61.120000 9.785000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 61.530000 9.785000 61.850000 ;
      LAYER met4 ;
        RECT 9.465000 61.530000 9.785000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 61.940000 9.785000 62.260000 ;
      LAYER met4 ;
        RECT 9.465000 61.940000 9.785000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 62.350000 9.785000 62.670000 ;
      LAYER met4 ;
        RECT 9.465000 62.350000 9.785000 62.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 58.250000 10.190000 58.570000 ;
      LAYER met4 ;
        RECT 9.870000 58.250000 10.190000 58.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 58.660000 10.190000 58.980000 ;
      LAYER met4 ;
        RECT 9.870000 58.660000 10.190000 58.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 59.070000 10.190000 59.390000 ;
      LAYER met4 ;
        RECT 9.870000 59.070000 10.190000 59.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 59.480000 10.190000 59.800000 ;
      LAYER met4 ;
        RECT 9.870000 59.480000 10.190000 59.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 59.890000 10.190000 60.210000 ;
      LAYER met4 ;
        RECT 9.870000 59.890000 10.190000 60.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 60.300000 10.190000 60.620000 ;
      LAYER met4 ;
        RECT 9.870000 60.300000 10.190000 60.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 60.710000 10.190000 61.030000 ;
      LAYER met4 ;
        RECT 9.870000 60.710000 10.190000 61.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 61.120000 10.190000 61.440000 ;
      LAYER met4 ;
        RECT 9.870000 61.120000 10.190000 61.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 61.530000 10.190000 61.850000 ;
      LAYER met4 ;
        RECT 9.870000 61.530000 10.190000 61.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 61.940000 10.190000 62.260000 ;
      LAYER met4 ;
        RECT 9.870000 61.940000 10.190000 62.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 62.350000 10.190000 62.670000 ;
      LAYER met4 ;
        RECT 9.870000 62.350000 10.190000 62.670000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.495000 25.840000 74.290000 200.000000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT 0.000000  2.135000 72.130000  15.035000 ;
      RECT 0.000000 15.035000 72.435000  19.885000 ;
      RECT 0.000000 19.885000 75.000000  30.385000 ;
      RECT 0.000000 30.385000 72.130000  36.835000 ;
      RECT 0.000000 36.835000 75.000000  40.085000 ;
      RECT 0.000000 40.085000 72.130000  58.335000 ;
      RECT 0.000000 58.335000 75.000000  62.585000 ;
      RECT 0.000000 62.585000 72.130000  96.585000 ;
      RECT 0.000000 96.585000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vssio_hvc
END LIBRARY
