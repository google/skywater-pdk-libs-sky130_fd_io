/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_SIO_MACRO_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_SIO_MACRO_PP_BLACKBOX_V

/**
 * top_sio_macro: sky130_fd_io__sio_macro consists of two SIO cells
 *                and a reference generator cell.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_sio_macro (
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           VINREF_DFT      ,
           VOUTREF_DFT     ,
           DFT_REFGEN      ,
           HLD_H_N_REFGEN  ,
           IBUF_SEL_REFGEN ,
           ENABLE_VDDA_H   ,
           ENABLE_H        ,
           VOHREF          ,
           VREG_EN_REFGEN  ,
           VTRIP_SEL_REFGEN,
           TIE_LO_ESD      ,
           IN_H            ,
           IN              ,
           PAD_A_NOESD_H   ,
           PAD             ,
           PAD_A_ESD_1_H   ,
           PAD_A_ESD_0_H   ,
           SLOW            ,
           VTRIP_SEL       ,
           HLD_H_N         ,
           VREG_EN         ,
           VOH_SEL         ,
           INP_DIS         ,
           HLD_OVR         ,
           OE_N            ,
           VREF_SEL        ,
           IBUF_SEL        ,
           DM0             ,
           DM1             ,
           OUT             ,
           VCCD            ,
           VCCHIB          ,
           VDDA            ,
           VDDIO           ,
           VDDIO_Q         ,
           VSSD            ,
           VSSIO           ,
           VSSIO_Q         ,
           VSWITCH         ,
           VSSA
       );

inout        AMUXBUS_A       ;
inout        AMUXBUS_B       ;
inout        VINREF_DFT      ;
inout        VOUTREF_DFT     ;
input        DFT_REFGEN      ;
input        HLD_H_N_REFGEN  ;
input        IBUF_SEL_REFGEN ;
input        ENABLE_VDDA_H   ;
input        ENABLE_H        ;
input        VOHREF          ;
input        VREG_EN_REFGEN  ;
input        VTRIP_SEL_REFGEN;
output [1:0] TIE_LO_ESD      ;
output [1:0] IN_H            ;
output [1:0] IN              ;
inout  [1:0] PAD_A_NOESD_H   ;
inout  [1:0] PAD             ;
inout  [1:0] PAD_A_ESD_1_H   ;
inout  [1:0] PAD_A_ESD_0_H   ;
input  [1:0] SLOW            ;
input  [1:0] VTRIP_SEL       ;
input  [1:0] HLD_H_N         ;
input  [1:0] VREG_EN         ;
input  [2:0] VOH_SEL         ;
input  [1:0] INP_DIS         ;
input  [1:0] HLD_OVR         ;
input  [1:0] OE_N            ;
input  [1:0] VREF_SEL        ;
input  [1:0] IBUF_SEL        ;
input  [2:0] DM0             ;
input  [2:0] DM1             ;
input  [1:0] OUT             ;
inout        VCCD            ;
inout        VCCHIB          ;
inout        VDDA            ;
inout        VDDIO           ;
inout        VDDIO_Q         ;
inout        VSSD            ;
inout        VSSIO           ;
inout        VSSIO_Q         ;
inout        VSWITCH         ;
inout        VSSA            ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_SIO_MACRO_PP_BLACKBOX_V
