# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_gpiov2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 80 BY 200 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430000 0.000000 62.690000 1.915000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865000  0.000000 46.195000 36.665000 ;
        RECT 45.865000 36.665000 46.195000 36.735000 ;
        RECT 45.865000 36.735000 46.265000 36.805000 ;
        RECT 45.965000 36.805000 46.335000 36.905000 ;
        RECT 46.065000 36.905000 46.435000 37.005000 ;
        RECT 46.070000 37.005000 46.535000 37.010000 ;
        RECT 46.220000 37.010000 48.225000 37.160000 ;
        RECT 46.370000 37.160000 48.075000 37.310000 ;
        RECT 46.400000 37.310000 48.045000 37.340000 ;
        RECT 47.910000 37.005000 48.375000 37.010000 ;
        RECT 47.960000 35.870000 48.740000 36.190000 ;
        RECT 47.975000 36.940000 48.380000 37.005000 ;
        RECT 48.040000 36.875000 48.445000 36.940000 ;
        RECT 48.070000 36.190000 48.630000 36.300000 ;
        RECT 48.110000 36.805000 48.510000 36.875000 ;
        RECT 48.180000 36.300000 48.520000 36.410000 ;
        RECT 48.180000 36.410000 48.515000 36.415000 ;
        RECT 48.180000 36.415000 48.510000 36.420000 ;
        RECT 48.180000 36.420000 48.510000 36.735000 ;
        RECT 48.180000 36.735000 48.510000 36.805000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.080000 57.360000 24.590000 57.430000 ;
        RECT 23.080000 57.430000 24.520000 57.500000 ;
        RECT 23.080000 57.500000 24.450000 57.570000 ;
        RECT 23.080000 57.570000 24.380000 57.640000 ;
        RECT 24.285000 57.345000 24.660000 57.360000 ;
        RECT 24.355000 57.275000 24.675000 57.345000 ;
        RECT 24.425000 57.205000 24.745000 57.275000 ;
        RECT 24.495000 57.135000 24.815000 57.205000 ;
        RECT 24.565000 57.065000 24.885000 57.135000 ;
        RECT 24.620000 57.010000 24.955000 57.065000 ;
        RECT 24.675000 53.255000 25.010000 53.310000 ;
        RECT 24.675000 53.310000 24.955000 53.365000 ;
        RECT 24.675000 53.365000 24.955000 56.955000 ;
        RECT 24.675000 56.955000 24.955000 57.010000 ;
        RECT 24.740000 53.190000 25.065000 53.255000 ;
        RECT 24.810000 53.120000 25.130000 53.190000 ;
        RECT 24.880000 53.050000 25.200000 53.120000 ;
        RECT 24.950000 52.980000 25.270000 53.050000 ;
        RECT 25.020000 52.910000 25.340000 52.980000 ;
        RECT 25.090000 52.840000 25.410000 52.910000 ;
        RECT 25.160000 52.770000 25.480000 52.840000 ;
        RECT 25.230000 52.700000 25.550000 52.770000 ;
        RECT 25.300000 52.630000 25.620000 52.700000 ;
        RECT 25.370000 52.560000 25.690000 52.630000 ;
        RECT 25.440000 52.490000 25.760000 52.560000 ;
        RECT 25.510000 52.420000 25.830000 52.490000 ;
        RECT 25.580000 52.350000 25.900000 52.420000 ;
        RECT 25.650000 52.280000 25.970000 52.350000 ;
        RECT 25.720000 52.210000 26.040000 52.280000 ;
        RECT 25.790000 52.140000 29.735000 52.210000 ;
        RECT 25.860000 52.070000 29.805000 52.140000 ;
        RECT 25.930000 52.000000 29.875000 52.070000 ;
        RECT 26.000000 51.930000 29.945000 52.000000 ;
        RECT 29.645000 51.910000 30.015000 51.930000 ;
        RECT 29.715000 51.840000 30.035000 51.910000 ;
        RECT 29.785000 51.770000 30.105000 51.840000 ;
        RECT 29.855000 51.700000 30.175000 51.770000 ;
        RECT 29.925000 51.630000 30.245000 51.700000 ;
        RECT 29.995000 51.560000 30.315000 51.630000 ;
        RECT 30.060000 51.495000 30.385000 51.560000 ;
        RECT 30.125000 17.630000 30.440000 17.685000 ;
        RECT 30.125000 17.685000 30.385000 17.740000 ;
        RECT 30.125000 17.740000 30.385000 36.345000 ;
        RECT 30.125000 36.345000 30.385000 36.400000 ;
        RECT 30.125000 36.400000 30.440000 36.455000 ;
        RECT 30.125000 38.010000 30.440000 38.065000 ;
        RECT 30.125000 38.065000 30.385000 38.120000 ;
        RECT 30.125000 38.120000 30.385000 51.430000 ;
        RECT 30.125000 51.430000 30.385000 51.495000 ;
        RECT 30.140000 37.995000 30.495000 38.010000 ;
        RECT 30.180000 17.575000 30.495000 17.630000 ;
        RECT 30.195000 36.455000 30.495000 36.525000 ;
        RECT 30.210000 37.925000 30.510000 37.995000 ;
        RECT 30.250000 17.505000 30.550000 17.575000 ;
        RECT 30.265000 36.525000 30.565000 36.595000 ;
        RECT 30.280000 36.595000 30.635000 36.610000 ;
        RECT 30.280000 37.855000 30.580000 37.925000 ;
        RECT 30.320000 17.435000 30.620000 17.505000 ;
        RECT 30.335000 36.610000 30.650000 36.665000 ;
        RECT 30.335000 37.800000 30.650000 37.855000 ;
        RECT 30.390000 17.365000 30.690000 17.435000 ;
        RECT 30.390000 36.665000 30.650000 36.720000 ;
        RECT 30.390000 36.720000 30.650000 37.745000 ;
        RECT 30.390000 37.745000 30.650000 37.800000 ;
        RECT 30.460000 17.295000 30.760000 17.365000 ;
        RECT 30.530000 17.225000 30.830000 17.295000 ;
        RECT 30.600000 17.155000 30.900000 17.225000 ;
        RECT 30.670000 17.085000 30.970000 17.155000 ;
        RECT 30.740000 17.015000 31.040000 17.085000 ;
        RECT 30.750000  0.000000 31.010000  2.155000 ;
        RECT 30.750000  2.155000 31.010000  2.210000 ;
        RECT 30.750000  2.210000 31.065000  2.265000 ;
        RECT 30.810000 16.945000 31.110000 17.015000 ;
        RECT 30.820000  2.265000 31.120000  2.335000 ;
        RECT 30.880000 16.875000 31.180000 16.945000 ;
        RECT 30.890000  2.335000 31.190000  2.405000 ;
        RECT 30.950000 16.805000 31.250000 16.875000 ;
        RECT 30.960000  2.405000 31.260000  2.475000 ;
        RECT 31.020000 16.735000 31.320000 16.805000 ;
        RECT 31.030000  2.475000 31.330000  2.545000 ;
        RECT 31.090000 16.665000 31.390000 16.735000 ;
        RECT 31.100000  2.545000 31.400000  2.615000 ;
        RECT 31.160000 16.595000 31.460000 16.665000 ;
        RECT 31.170000  2.615000 31.470000  2.685000 ;
        RECT 31.195000  2.685000 31.540000  2.710000 ;
        RECT 31.230000 16.525000 31.530000 16.595000 ;
        RECT 31.250000  2.710000 31.565000  2.765000 ;
        RECT 31.300000 16.455000 31.600000 16.525000 ;
        RECT 31.305000  2.765000 31.565000  2.820000 ;
        RECT 31.305000  2.820000 31.565000  4.335000 ;
        RECT 31.305000  4.335000 31.565000  4.390000 ;
        RECT 31.305000  4.390000 31.620000  4.445000 ;
        RECT 31.370000 16.385000 31.670000 16.455000 ;
        RECT 31.375000  4.445000 31.675000  4.515000 ;
        RECT 31.440000 16.315000 31.740000 16.385000 ;
        RECT 31.445000  4.515000 31.745000  4.585000 ;
        RECT 31.510000 16.245000 31.810000 16.315000 ;
        RECT 31.515000  4.585000 31.815000  4.655000 ;
        RECT 31.580000  4.655000 31.885000  4.720000 ;
        RECT 31.580000 16.175000 31.880000 16.245000 ;
        RECT 31.635000  4.720000 31.950000  4.775000 ;
        RECT 31.635000 16.120000 31.950000 16.175000 ;
        RECT 31.690000  4.775000 31.950000  4.830000 ;
        RECT 31.690000  4.830000 31.950000 16.065000 ;
        RECT 31.690000 16.065000 31.950000 16.120000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.590000 0.545000 50.360000 0.825000 ;
        RECT 49.625000 0.510000 50.325000 0.545000 ;
        RECT 49.695000 0.440000 50.255000 0.510000 ;
        RECT 49.765000 0.370000 50.185000 0.440000 ;
        RECT 49.835000 0.300000 50.115000 0.370000 ;
        RECT 49.845000 0.290000 50.115000 0.300000 ;
        RECT 49.855000 0.000000 50.115000 0.280000 ;
        RECT 49.855000 0.280000 50.115000 0.290000 ;
    END
  END DM[0]
  PIN DM[1]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.540000 1.195000 67.360000 1.475000 ;
        RECT 66.595000 1.140000 67.305000 1.195000 ;
        RECT 66.665000 1.070000 67.235000 1.140000 ;
        RECT 66.735000 1.000000 67.165000 1.070000 ;
        RECT 66.805000 0.930000 67.095000 1.000000 ;
        RECT 66.820000 0.915000 67.095000 0.930000 ;
        RECT 66.835000 0.000000 67.095000 0.900000 ;
        RECT 66.835000 0.900000 67.095000 0.915000 ;
    END
  END DM[1]
  PIN DM[2]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490000 0.000000 28.750000 3.960000 ;
        RECT 28.490000 3.960000 28.750000 4.015000 ;
        RECT 28.490000 4.015000 28.805000 4.070000 ;
        RECT 28.560000 4.070000 28.860000 4.140000 ;
        RECT 28.630000 4.140000 28.930000 4.210000 ;
        RECT 28.700000 4.210000 29.000000 4.280000 ;
        RECT 28.770000 4.280000 29.070000 4.350000 ;
        RECT 28.840000 4.350000 29.140000 4.420000 ;
        RECT 28.910000 4.420000 29.210000 4.490000 ;
        RECT 28.980000 4.490000 29.280000 4.560000 ;
        RECT 29.050000 4.560000 29.350000 4.630000 ;
        RECT 29.100000 4.630000 29.420000 4.680000 ;
        RECT 29.155000 4.680000 29.470000 4.735000 ;
        RECT 29.210000 4.735000 29.470000 4.790000 ;
        RECT 29.210000 4.790000 29.470000 6.780000 ;
    END
  END DM[2]
  PIN ENABLE_H
    ANTENNAGATEAREA  4.860000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.135000 2.225000 35.450000 2.280000 ;
        RECT 35.135000 2.280000 35.395000 2.335000 ;
        RECT 35.135000 2.335000 35.395000 3.885000 ;
        RECT 35.140000 2.220000 35.505000 2.225000 ;
        RECT 35.210000 2.150000 35.510000 2.220000 ;
        RECT 35.280000 2.080000 35.580000 2.150000 ;
        RECT 35.350000 2.010000 35.650000 2.080000 ;
        RECT 35.405000 1.955000 35.720000 2.010000 ;
        RECT 35.460000 0.000000 35.720000 1.900000 ;
        RECT 35.460000 1.900000 35.720000 1.955000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390000 0.000000 38.650000 3.715000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  3.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.315000 56.460000  7.630000 56.515000 ;
        RECT  7.315000 56.515000  7.575000 56.570000 ;
        RECT  7.315000 56.570000  7.575000 73.615000 ;
        RECT  7.315000 73.615000  7.575000 73.670000 ;
        RECT  7.315000 73.670000  7.630000 73.725000 ;
        RECT  7.375000 56.400000  7.685000 56.460000 ;
        RECT  7.385000 73.725000  7.685000 73.795000 ;
        RECT  7.445000 56.330000  7.745000 56.400000 ;
        RECT  7.455000 73.795000  7.755000 73.865000 ;
        RECT  7.515000 56.260000  7.815000 56.330000 ;
        RECT  7.525000 73.865000  7.825000 73.935000 ;
        RECT  7.585000 56.190000  7.885000 56.260000 ;
        RECT  7.595000 73.935000  7.895000 74.005000 ;
        RECT  7.655000 56.120000  7.955000 56.190000 ;
        RECT  7.665000 74.005000  7.965000 74.075000 ;
        RECT  7.695000 74.075000  8.035000 74.105000 ;
        RECT  7.725000 56.050000  8.025000 56.120000 ;
        RECT  7.750000 74.105000  8.065000 74.160000 ;
        RECT  7.795000 55.980000  8.095000 56.050000 ;
        RECT  7.805000 74.160000  8.065000 74.215000 ;
        RECT  7.805000 74.215000  8.065000 74.680000 ;
        RECT  7.805000 74.680000  8.065000 74.735000 ;
        RECT  7.805000 74.735000  8.120000 74.790000 ;
        RECT  7.865000 55.910000  8.165000 55.980000 ;
        RECT  7.875000 74.790000  8.175000 74.860000 ;
        RECT  7.920000 55.855000  8.235000 55.910000 ;
        RECT  7.920000 77.285000  8.560000 77.545000 ;
        RECT  7.945000 74.860000  8.245000 74.930000 ;
        RECT  7.975000 53.960000  8.290000 54.015000 ;
        RECT  7.975000 54.015000  8.235000 54.070000 ;
        RECT  7.975000 54.070000  8.235000 55.800000 ;
        RECT  7.975000 55.800000  8.235000 55.855000 ;
        RECT  8.015000 74.930000  8.315000 75.000000 ;
        RECT  8.030000 53.905000  8.345000 53.960000 ;
        RECT  8.085000 53.850000  8.400000 53.905000 ;
        RECT  8.085000 75.000000  8.385000 75.070000 ;
        RECT  8.085000 77.240000  8.515000 77.285000 ;
        RECT  8.100000 75.070000  8.455000 75.085000 ;
        RECT  8.130000 77.195000  8.470000 77.240000 ;
        RECT  8.140000 53.795000  8.455000 53.850000 ;
        RECT  8.155000 75.085000  8.470000 75.140000 ;
        RECT  8.170000 77.155000  8.470000 77.195000 ;
        RECT  8.195000 44.075000  8.510000 44.130000 ;
        RECT  8.195000 44.130000  8.455000 44.185000 ;
        RECT  8.195000 44.185000  8.455000 53.740000 ;
        RECT  8.195000 53.740000  8.455000 53.795000 ;
        RECT  8.210000 44.060000  8.565000 44.075000 ;
        RECT  8.210000 75.140000  8.470000 75.195000 ;
        RECT  8.210000 75.195000  8.470000 77.115000 ;
        RECT  8.210000 77.115000  8.470000 77.155000 ;
        RECT  8.280000 43.990000  8.580000 44.060000 ;
        RECT  8.350000 43.920000  8.650000 43.990000 ;
        RECT  8.420000 43.850000  8.720000 43.920000 ;
        RECT  8.490000 43.780000  8.790000 43.850000 ;
        RECT  8.560000 43.710000  8.860000 43.780000 ;
        RECT  8.630000 43.640000  8.930000 43.710000 ;
        RECT  8.700000 43.570000  9.000000 43.640000 ;
        RECT  8.770000 43.500000  9.070000 43.570000 ;
        RECT  8.840000 43.430000  9.140000 43.500000 ;
        RECT  8.910000 43.360000  9.210000 43.430000 ;
        RECT  8.980000 43.290000  9.280000 43.360000 ;
        RECT  9.050000 43.220000  9.350000 43.290000 ;
        RECT  9.120000 43.150000  9.420000 43.220000 ;
        RECT  9.190000 43.080000  9.490000 43.150000 ;
        RECT  9.260000 43.010000  9.560000 43.080000 ;
        RECT  9.330000 42.940000  9.630000 43.010000 ;
        RECT  9.400000 42.870000  9.700000 42.940000 ;
        RECT  9.470000 42.800000  9.770000 42.870000 ;
        RECT  9.540000 42.730000  9.840000 42.800000 ;
        RECT  9.610000 42.660000  9.910000 42.730000 ;
        RECT  9.680000 42.590000  9.980000 42.660000 ;
        RECT  9.750000 42.520000 10.050000 42.590000 ;
        RECT  9.820000 42.450000 10.120000 42.520000 ;
        RECT  9.890000 42.380000 10.190000 42.450000 ;
        RECT  9.960000 42.310000 10.260000 42.380000 ;
        RECT 10.030000 42.240000 10.330000 42.310000 ;
        RECT 10.100000 42.170000 10.400000 42.240000 ;
        RECT 10.170000 42.100000 10.470000 42.170000 ;
        RECT 10.240000 42.030000 10.540000 42.100000 ;
        RECT 10.310000 41.960000 10.610000 42.030000 ;
        RECT 10.380000 41.890000 10.680000 41.960000 ;
        RECT 10.450000 41.820000 10.750000 41.890000 ;
        RECT 10.520000 41.750000 10.820000 41.820000 ;
        RECT 10.590000 41.680000 10.890000 41.750000 ;
        RECT 10.660000 41.610000 10.960000 41.680000 ;
        RECT 10.730000 41.540000 11.030000 41.610000 ;
        RECT 10.800000 41.470000 11.100000 41.540000 ;
        RECT 10.870000 41.400000 11.170000 41.470000 ;
        RECT 10.940000 41.330000 11.240000 41.400000 ;
        RECT 11.010000 41.260000 11.310000 41.330000 ;
        RECT 11.080000 41.190000 11.380000 41.260000 ;
        RECT 11.150000 41.120000 11.450000 41.190000 ;
        RECT 11.220000 41.050000 11.520000 41.120000 ;
        RECT 11.290000 40.980000 11.590000 41.050000 ;
        RECT 11.360000 40.910000 11.660000 40.980000 ;
        RECT 11.430000 40.840000 11.730000 40.910000 ;
        RECT 11.500000 40.770000 11.800000 40.840000 ;
        RECT 11.570000 40.700000 11.870000 40.770000 ;
        RECT 11.640000 40.630000 11.940000 40.700000 ;
        RECT 11.710000 40.560000 12.010000 40.630000 ;
        RECT 11.780000 40.490000 12.080000 40.560000 ;
        RECT 11.850000 40.420000 12.150000 40.490000 ;
        RECT 11.920000 40.350000 12.220000 40.420000 ;
        RECT 11.990000 40.280000 12.290000 40.350000 ;
        RECT 12.060000 40.210000 12.360000 40.280000 ;
        RECT 12.130000 40.140000 12.430000 40.210000 ;
        RECT 12.200000 40.070000 12.500000 40.140000 ;
        RECT 12.270000 40.000000 12.570000 40.070000 ;
        RECT 12.340000 39.930000 12.640000 40.000000 ;
        RECT 12.410000 39.860000 12.710000 39.930000 ;
        RECT 12.480000 39.790000 12.780000 39.860000 ;
        RECT 12.550000 39.720000 12.850000 39.790000 ;
        RECT 12.620000 39.650000 12.920000 39.720000 ;
        RECT 12.690000 39.580000 12.990000 39.650000 ;
        RECT 12.755000  0.000000 13.015000  5.240000 ;
        RECT 12.755000  5.240000 13.015000  5.295000 ;
        RECT 12.755000  5.295000 13.070000  5.350000 ;
        RECT 12.760000 39.510000 13.060000 39.580000 ;
        RECT 12.825000  5.350000 13.125000  5.420000 ;
        RECT 12.830000 39.440000 13.130000 39.510000 ;
        RECT 12.895000  5.420000 13.195000  5.490000 ;
        RECT 12.900000 39.370000 13.200000 39.440000 ;
        RECT 12.965000  5.490000 13.265000  5.560000 ;
        RECT 12.970000 39.300000 13.270000 39.370000 ;
        RECT 13.035000  5.560000 13.335000  5.630000 ;
        RECT 13.040000 39.230000 13.340000 39.300000 ;
        RECT 13.105000  5.630000 13.405000  5.700000 ;
        RECT 13.110000 39.160000 13.410000 39.230000 ;
        RECT 13.175000  5.700000 13.475000  5.770000 ;
        RECT 13.180000 39.090000 13.480000 39.160000 ;
        RECT 13.245000  5.770000 13.545000  5.840000 ;
        RECT 13.250000 39.020000 13.550000 39.090000 ;
        RECT 13.315000  5.840000 13.615000  5.910000 ;
        RECT 13.320000 38.950000 13.620000 39.020000 ;
        RECT 13.385000  5.910000 13.685000  5.980000 ;
        RECT 13.390000 38.880000 13.690000 38.950000 ;
        RECT 13.455000  5.980000 13.755000  6.050000 ;
        RECT 13.460000 38.810000 13.760000 38.880000 ;
        RECT 13.525000  6.050000 13.825000  6.120000 ;
        RECT 13.530000 38.740000 13.830000 38.810000 ;
        RECT 13.595000  6.120000 13.895000  6.190000 ;
        RECT 13.600000 38.670000 13.900000 38.740000 ;
        RECT 13.665000  6.190000 13.965000  6.260000 ;
        RECT 13.670000 38.600000 13.970000 38.670000 ;
        RECT 13.735000  6.260000 14.035000  6.330000 ;
        RECT 13.740000 38.530000 14.040000 38.600000 ;
        RECT 13.805000  6.330000 14.105000  6.400000 ;
        RECT 13.810000 38.460000 14.110000 38.530000 ;
        RECT 13.860000  6.400000 14.175000  6.455000 ;
        RECT 13.880000 38.390000 14.180000 38.460000 ;
        RECT 13.915000  6.455000 14.230000  6.510000 ;
        RECT 13.950000 38.320000 14.250000 38.390000 ;
        RECT 13.970000  6.510000 14.230000  6.565000 ;
        RECT 13.970000  6.565000 14.230000 18.115000 ;
        RECT 13.970000 18.115000 14.230000 18.170000 ;
        RECT 13.970000 18.170000 14.285000 18.225000 ;
        RECT 14.020000 38.250000 14.320000 38.320000 ;
        RECT 14.040000 18.225000 14.340000 18.295000 ;
        RECT 14.090000 38.180000 14.390000 38.250000 ;
        RECT 14.110000 18.295000 14.410000 18.365000 ;
        RECT 14.160000 38.110000 14.460000 38.180000 ;
        RECT 14.180000 18.365000 14.480000 18.435000 ;
        RECT 14.230000 38.040000 14.530000 38.110000 ;
        RECT 14.250000 18.435000 14.550000 18.505000 ;
        RECT 14.300000 37.970000 14.600000 38.040000 ;
        RECT 14.320000 18.505000 14.620000 18.575000 ;
        RECT 14.370000 37.900000 14.670000 37.970000 ;
        RECT 14.390000 18.575000 14.690000 18.645000 ;
        RECT 14.440000 37.830000 14.740000 37.900000 ;
        RECT 14.460000 18.645000 14.760000 18.715000 ;
        RECT 14.510000 37.760000 14.810000 37.830000 ;
        RECT 14.530000 18.715000 14.830000 18.785000 ;
        RECT 14.580000 37.690000 14.880000 37.760000 ;
        RECT 14.600000 18.785000 14.900000 18.855000 ;
        RECT 14.650000 37.620000 14.950000 37.690000 ;
        RECT 14.670000 18.855000 14.970000 18.925000 ;
        RECT 14.720000 37.550000 15.020000 37.620000 ;
        RECT 14.740000 18.925000 15.040000 18.995000 ;
        RECT 14.790000 37.480000 15.090000 37.550000 ;
        RECT 14.810000 18.995000 15.110000 19.065000 ;
        RECT 14.860000 37.410000 15.160000 37.480000 ;
        RECT 14.880000 19.065000 15.180000 19.135000 ;
        RECT 14.915000 37.355000 15.230000 37.410000 ;
        RECT 14.950000 19.135000 15.250000 19.205000 ;
        RECT 14.970000 31.960000 15.285000 32.015000 ;
        RECT 14.970000 32.015000 15.230000 32.070000 ;
        RECT 14.970000 32.070000 15.230000 37.300000 ;
        RECT 14.970000 37.300000 15.230000 37.355000 ;
        RECT 14.995000 31.935000 15.340000 31.960000 ;
        RECT 15.020000 19.205000 15.320000 19.275000 ;
        RECT 15.065000 31.865000 15.365000 31.935000 ;
        RECT 15.090000 19.275000 15.390000 19.345000 ;
        RECT 15.135000 31.795000 15.435000 31.865000 ;
        RECT 15.160000 19.345000 15.460000 19.415000 ;
        RECT 15.205000 31.725000 15.505000 31.795000 ;
        RECT 15.230000 19.415000 15.530000 19.485000 ;
        RECT 15.275000 19.485000 15.600000 19.530000 ;
        RECT 15.275000 31.655000 15.575000 31.725000 ;
        RECT 15.330000 19.530000 15.645000 19.585000 ;
        RECT 15.330000 31.600000 15.645000 31.655000 ;
        RECT 15.385000 19.585000 15.645000 19.640000 ;
        RECT 15.385000 19.640000 15.645000 31.545000 ;
        RECT 15.385000 31.545000 15.645000 31.600000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580000 0.000000 78.910000 176.480000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    ANTENNAGATEAREA  3.120000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.250000 43.835000 11.565000 43.890000 ;
        RECT 11.250000 43.890000 11.510000 43.945000 ;
        RECT 11.250000 43.945000 11.510000 47.275000 ;
        RECT 11.250000 47.275000 11.510000 47.330000 ;
        RECT 11.250000 47.330000 11.565000 47.385000 ;
        RECT 11.270000 43.815000 11.620000 43.835000 ;
        RECT 11.320000 47.385000 11.620000 47.455000 ;
        RECT 11.340000 43.745000 11.640000 43.815000 ;
        RECT 11.390000 47.455000 11.690000 47.525000 ;
        RECT 11.410000 43.675000 11.710000 43.745000 ;
        RECT 11.460000 47.525000 11.760000 47.595000 ;
        RECT 11.480000 43.605000 11.780000 43.675000 ;
        RECT 11.530000 47.595000 11.830000 47.665000 ;
        RECT 11.550000 43.535000 11.850000 43.605000 ;
        RECT 11.600000 47.665000 11.900000 47.735000 ;
        RECT 11.620000 43.465000 11.920000 43.535000 ;
        RECT 11.670000 47.735000 11.970000 47.805000 ;
        RECT 11.680000 47.805000 12.040000 47.815000 ;
        RECT 11.690000 43.395000 11.990000 43.465000 ;
        RECT 11.750000 47.815000 13.850000 47.885000 ;
        RECT 11.760000 43.325000 12.060000 43.395000 ;
        RECT 11.820000 47.885000 13.920000 47.955000 ;
        RECT 11.830000 43.255000 12.130000 43.325000 ;
        RECT 11.890000 47.955000 13.990000 48.025000 ;
        RECT 11.900000 43.185000 12.200000 43.255000 ;
        RECT 11.940000 48.025000 14.060000 48.075000 ;
        RECT 11.970000 43.115000 12.270000 43.185000 ;
        RECT 12.040000 43.045000 12.340000 43.115000 ;
        RECT 12.110000 42.975000 12.410000 43.045000 ;
        RECT 12.180000 42.905000 12.480000 42.975000 ;
        RECT 12.250000 42.835000 12.550000 42.905000 ;
        RECT 12.320000 42.765000 12.620000 42.835000 ;
        RECT 12.390000 42.695000 12.690000 42.765000 ;
        RECT 12.460000 42.625000 12.760000 42.695000 ;
        RECT 12.530000 42.555000 12.830000 42.625000 ;
        RECT 12.600000 42.485000 12.900000 42.555000 ;
        RECT 12.670000 42.415000 12.970000 42.485000 ;
        RECT 12.740000 42.345000 13.040000 42.415000 ;
        RECT 12.810000 42.275000 13.110000 42.345000 ;
        RECT 12.880000 42.205000 13.180000 42.275000 ;
        RECT 12.950000 42.135000 13.250000 42.205000 ;
        RECT 13.020000 42.065000 13.320000 42.135000 ;
        RECT 13.090000 41.995000 13.390000 42.065000 ;
        RECT 13.160000 41.925000 13.460000 41.995000 ;
        RECT 13.230000 41.855000 13.530000 41.925000 ;
        RECT 13.300000 41.785000 13.600000 41.855000 ;
        RECT 13.370000 41.715000 13.670000 41.785000 ;
        RECT 13.440000 41.645000 13.740000 41.715000 ;
        RECT 13.510000 41.575000 13.810000 41.645000 ;
        RECT 13.565000 41.520000 13.880000 41.575000 ;
        RECT 13.620000 40.430000 13.935000 40.485000 ;
        RECT 13.620000 40.485000 13.880000 40.540000 ;
        RECT 13.620000 40.540000 13.880000 41.465000 ;
        RECT 13.620000 41.465000 13.880000 41.520000 ;
        RECT 13.640000 40.410000 13.990000 40.430000 ;
        RECT 13.710000 40.340000 14.010000 40.410000 ;
        RECT 13.780000 40.270000 14.080000 40.340000 ;
        RECT 13.810000 48.075000 14.110000 48.145000 ;
        RECT 13.850000 40.200000 14.150000 40.270000 ;
        RECT 13.880000 48.145000 14.180000 48.215000 ;
        RECT 13.920000 40.130000 14.220000 40.200000 ;
        RECT 13.950000 48.215000 14.250000 48.285000 ;
        RECT 13.990000 40.060000 14.290000 40.130000 ;
        RECT 14.020000 48.285000 14.320000 48.355000 ;
        RECT 14.060000 39.990000 14.360000 40.060000 ;
        RECT 14.090000 48.355000 14.390000 48.425000 ;
        RECT 14.130000 39.920000 14.430000 39.990000 ;
        RECT 14.160000 48.425000 14.460000 48.495000 ;
        RECT 14.180000 39.870000 15.420000 39.920000 ;
        RECT 14.195000 58.050000 14.835000 58.310000 ;
        RECT 14.210000 58.035000 14.820000 58.050000 ;
        RECT 14.230000 48.495000 14.530000 48.565000 ;
        RECT 14.240000 48.565000 14.600000 48.575000 ;
        RECT 14.250000 39.800000 15.470000 39.870000 ;
        RECT 14.280000 57.965000 14.750000 58.035000 ;
        RECT 14.295000 48.575000 14.610000 48.630000 ;
        RECT 14.320000 39.730000 15.540000 39.800000 ;
        RECT 14.350000 48.630000 14.610000 48.685000 ;
        RECT 14.350000 48.685000 14.610000 57.825000 ;
        RECT 14.350000 57.825000 14.610000 57.860000 ;
        RECT 14.350000 57.860000 14.645000 57.895000 ;
        RECT 14.350000 57.895000 14.680000 57.965000 ;
        RECT 14.390000 39.660000 15.610000 39.730000 ;
        RECT 15.365000 39.605000 15.680000 39.660000 ;
        RECT 15.435000 39.535000 15.735000 39.605000 ;
        RECT 15.505000 39.465000 15.805000 39.535000 ;
        RECT 15.575000 39.395000 15.875000 39.465000 ;
        RECT 15.645000 39.325000 15.945000 39.395000 ;
        RECT 15.715000 39.255000 16.015000 39.325000 ;
        RECT 15.785000 39.185000 16.085000 39.255000 ;
        RECT 15.855000 39.115000 16.155000 39.185000 ;
        RECT 15.925000 39.045000 16.225000 39.115000 ;
        RECT 15.995000 38.975000 16.295000 39.045000 ;
        RECT 16.065000 38.905000 16.365000 38.975000 ;
        RECT 16.135000 38.835000 16.435000 38.905000 ;
        RECT 16.205000 38.765000 16.505000 38.835000 ;
        RECT 16.275000 38.695000 16.575000 38.765000 ;
        RECT 16.310000  0.000000 16.570000  2.210000 ;
        RECT 16.310000  2.210000 16.570000  2.265000 ;
        RECT 16.310000  2.265000 16.625000  2.320000 ;
        RECT 16.345000 38.625000 16.645000 38.695000 ;
        RECT 16.365000 31.560000 16.680000 31.615000 ;
        RECT 16.365000 31.615000 16.625000 31.670000 ;
        RECT 16.365000 31.670000 16.625000 34.210000 ;
        RECT 16.365000 34.210000 16.625000 34.265000 ;
        RECT 16.365000 34.265000 16.680000 34.320000 ;
        RECT 16.370000 31.555000 16.735000 31.560000 ;
        RECT 16.380000  2.320000 16.680000  2.390000 ;
        RECT 16.415000 38.555000 16.715000 38.625000 ;
        RECT 16.435000 31.490000 16.740000 31.555000 ;
        RECT 16.435000 34.320000 16.735000 34.390000 ;
        RECT 16.450000  2.390000 16.750000  2.460000 ;
        RECT 16.485000 38.485000 16.785000 38.555000 ;
        RECT 16.500000 31.425000 16.805000 31.490000 ;
        RECT 16.505000 34.390000 16.805000 34.460000 ;
        RECT 16.520000  2.460000 16.820000  2.530000 ;
        RECT 16.555000 31.370000 16.870000 31.425000 ;
        RECT 16.555000 38.415000 16.855000 38.485000 ;
        RECT 16.575000 34.460000 16.875000 34.530000 ;
        RECT 16.590000  2.530000 16.890000  2.600000 ;
        RECT 16.610000  7.160000 16.925000  7.215000 ;
        RECT 16.610000  7.215000 16.870000  7.270000 ;
        RECT 16.610000  7.270000 16.870000 11.540000 ;
        RECT 16.610000 12.475000 16.870000 31.315000 ;
        RECT 16.610000 31.315000 16.870000 31.370000 ;
        RECT 16.615000 12.470000 16.870000 12.475000 ;
        RECT 16.625000 38.345000 16.925000 38.415000 ;
        RECT 16.635000  7.135000 16.980000  7.160000 ;
        RECT 16.645000 34.530000 16.945000 34.600000 ;
        RECT 16.655000 11.540000 16.870000 11.585000 ;
        RECT 16.660000  2.600000 16.960000  2.670000 ;
        RECT 16.660000 12.425000 16.870000 12.470000 ;
        RECT 16.695000 38.275000 16.995000 38.345000 ;
        RECT 16.700000 11.585000 16.870000 11.630000 ;
        RECT 16.705000  7.065000 17.005000  7.135000 ;
        RECT 16.705000 11.630000 16.870000 11.635000 ;
        RECT 16.705000 11.635000 16.870000 12.380000 ;
        RECT 16.705000 12.380000 16.870000 12.425000 ;
        RECT 16.715000 34.600000 17.015000 34.670000 ;
        RECT 16.730000  2.670000 17.030000  2.740000 ;
        RECT 16.765000 38.205000 17.065000 38.275000 ;
        RECT 16.775000  6.995000 17.075000  7.065000 ;
        RECT 16.785000 34.670000 17.085000 34.740000 ;
        RECT 16.800000  2.740000 17.100000  2.810000 ;
        RECT 16.835000 38.135000 17.135000 38.205000 ;
        RECT 16.845000  6.925000 17.145000  6.995000 ;
        RECT 16.855000 34.740000 17.155000 34.810000 ;
        RECT 16.870000  2.810000 17.170000  2.880000 ;
        RECT 16.905000 38.065000 17.205000 38.135000 ;
        RECT 16.915000  6.855000 17.215000  6.925000 ;
        RECT 16.925000 34.810000 17.225000 34.880000 ;
        RECT 16.940000  2.880000 17.240000  2.950000 ;
        RECT 16.975000 37.995000 17.275000 38.065000 ;
        RECT 16.985000  2.950000 17.310000  2.995000 ;
        RECT 16.985000  6.785000 17.285000  6.855000 ;
        RECT 16.995000 34.880000 17.295000 34.950000 ;
        RECT 17.040000  2.995000 17.355000  3.050000 ;
        RECT 17.040000  6.730000 17.355000  6.785000 ;
        RECT 17.045000 37.925000 17.345000 37.995000 ;
        RECT 17.065000 34.950000 17.365000 35.020000 ;
        RECT 17.095000  3.050000 17.355000  3.105000 ;
        RECT 17.095000  3.105000 17.355000  6.675000 ;
        RECT 17.095000  6.675000 17.355000  6.730000 ;
        RECT 17.115000 37.855000 17.415000 37.925000 ;
        RECT 17.135000 35.020000 17.435000 35.090000 ;
        RECT 17.185000 37.785000 17.485000 37.855000 ;
        RECT 17.205000 35.090000 17.505000 35.160000 ;
        RECT 17.255000 37.715000 17.555000 37.785000 ;
        RECT 17.275000 35.160000 17.575000 35.230000 ;
        RECT 17.325000 37.645000 17.625000 37.715000 ;
        RECT 17.345000 35.230000 17.645000 35.300000 ;
        RECT 17.395000 37.575000 17.695000 37.645000 ;
        RECT 17.415000 35.300000 17.715000 35.370000 ;
        RECT 17.465000 35.370000 17.785000 35.420000 ;
        RECT 17.465000 37.505000 17.765000 37.575000 ;
        RECT 17.520000 35.420000 17.835000 35.475000 ;
        RECT 17.520000 37.450000 17.835000 37.505000 ;
        RECT 17.575000 35.475000 17.835000 35.530000 ;
        RECT 17.575000 35.530000 17.835000 37.395000 ;
        RECT 17.575000 37.395000 17.835000 37.450000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    ANTENNAGATEAREA  1.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815000 0.000000 32.075000 3.965000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600000 0.000000 26.860000 1.695000 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420000 0.000000 5.650000 4.375000 ;
        RECT 5.420000 4.375000 5.650000 4.425000 ;
        RECT 5.420000 4.425000 5.700000 4.475000 ;
        RECT 5.490000 4.475000 5.750000 4.545000 ;
        RECT 5.560000 4.545000 5.820000 4.615000 ;
        RECT 5.630000 4.615000 5.890000 4.685000 ;
        RECT 5.700000 4.685000 5.960000 4.755000 ;
        RECT 5.770000 4.755000 6.030000 4.825000 ;
        RECT 5.840000 4.825000 6.100000 4.895000 ;
        RECT 5.910000 4.895000 6.170000 4.965000 ;
        RECT 5.910000 6.425000 6.550000 6.685000 ;
        RECT 5.980000 4.965000 6.240000 5.035000 ;
        RECT 6.050000 5.035000 6.310000 5.105000 ;
        RECT 6.120000 5.105000 6.380000 5.175000 ;
        RECT 6.180000 6.390000 6.550000 6.425000 ;
        RECT 6.190000 5.175000 6.450000 5.245000 ;
        RECT 6.220000 5.245000 6.520000 5.275000 ;
        RECT 6.250000 6.320000 6.550000 6.390000 ;
        RECT 6.270000 5.275000 6.550000 5.325000 ;
        RECT 6.320000 5.325000 6.550000 5.375000 ;
        RECT 6.320000 5.375000 6.550000 6.250000 ;
        RECT 6.320000 6.250000 6.550000 6.320000 ;
    END
  END IB_MODE_SEL
  PIN IN
    ANTENNAPARTIALMETALSIDEAREA  303.1200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240000 0.000000 79.570000 176.480000 ;
    END
  END IN
  PIN INP_DIS
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245000 0.000000 45.505000 4.980000 ;
        RECT 45.245000 4.980000 45.505000 5.035000 ;
        RECT 45.245000 5.035000 45.560000 5.090000 ;
        RECT 45.315000 5.090000 45.615000 5.160000 ;
        RECT 45.385000 5.160000 45.685000 5.230000 ;
        RECT 45.455000 5.230000 45.755000 5.300000 ;
        RECT 45.525000 5.300000 45.825000 5.370000 ;
        RECT 45.595000 5.370000 45.895000 5.440000 ;
        RECT 45.665000 5.440000 45.965000 5.510000 ;
        RECT 45.735000 5.510000 46.035000 5.580000 ;
        RECT 45.745000 5.580000 46.105000 5.590000 ;
        RECT 45.800000 5.590000 46.115000 5.645000 ;
        RECT 45.855000 5.645000 46.115000 5.700000 ;
        RECT 45.855000 5.700000 46.115000 6.780000 ;
    END
  END INP_DIS
  PIN IN_H
    ANTENNAPARTIALMETALSIDEAREA  291.9480 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400000   0.000000 1.020000 178.235000 ;
        RECT 0.400000 178.235000 1.020000 178.360000 ;
        RECT 0.400000 178.360000 1.145000 178.485000 ;
        RECT 0.550000 178.485000 1.270000 178.635000 ;
        RECT 0.700000 178.635000 1.420000 178.785000 ;
        RECT 0.850000 178.785000 1.570000 178.935000 ;
        RECT 1.000000 178.935000 1.720000 179.085000 ;
        RECT 1.150000 179.085000 1.870000 179.235000 ;
        RECT 1.300000 179.235000 2.020000 179.385000 ;
        RECT 1.450000 179.385000 2.170000 179.535000 ;
        RECT 1.600000 179.535000 2.320000 179.685000 ;
        RECT 1.750000 179.685000 2.470000 179.835000 ;
        RECT 1.900000 179.835000 2.620000 179.985000 ;
        RECT 2.050000 179.985000 2.770000 180.135000 ;
        RECT 2.200000 180.135000 2.920000 180.285000 ;
        RECT 2.350000 180.285000 3.070000 180.435000 ;
        RECT 2.355000 180.435000 3.220000 180.440000 ;
        RECT 2.505000 180.440000 4.565000 180.590000 ;
        RECT 2.655000 180.590000 4.565000 180.740000 ;
        RECT 2.805000 180.740000 4.565000 180.890000 ;
        RECT 2.955000 180.890000 4.565000 181.040000 ;
        RECT 3.085000 181.040000 4.565000 181.170000 ;
    END
  END IN_H
  PIN OE_N
    ANTENNAGATEAREA  1.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375000  0.000000 3.605000  4.375000 ;
        RECT 3.375000  4.375000 3.605000  4.425000 ;
        RECT 3.375000  4.425000 3.655000  4.475000 ;
        RECT 3.445000  4.475000 3.705000  4.545000 ;
        RECT 3.515000  4.545000 3.775000  4.615000 ;
        RECT 3.585000  4.615000 3.845000  4.685000 ;
        RECT 3.655000  4.685000 3.915000  4.755000 ;
        RECT 3.725000  4.755000 3.985000  4.825000 ;
        RECT 3.770000  4.825000 4.055000  4.870000 ;
        RECT 3.840000  4.870000 5.225000  4.940000 ;
        RECT 3.910000  4.940000 5.295000  5.010000 ;
        RECT 3.980000  5.010000 5.365000  5.080000 ;
        RECT 4.000000  5.080000 5.435000  5.100000 ;
        RECT 5.195000  5.100000 5.455000  5.170000 ;
        RECT 5.265000  5.170000 5.525000  5.240000 ;
        RECT 5.300000  5.240000 5.595000  5.275000 ;
        RECT 5.350000  5.275000 5.630000  5.325000 ;
        RECT 5.400000  5.325000 5.630000  5.375000 ;
        RECT 5.400000  5.375000 5.630000  8.250000 ;
        RECT 5.400000  8.250000 5.630000  8.300000 ;
        RECT 5.400000  8.300000 5.680000  8.350000 ;
        RECT 5.470000  8.350000 5.730000  8.420000 ;
        RECT 5.540000  8.420000 5.800000  8.490000 ;
        RECT 5.610000  8.490000 5.870000  8.560000 ;
        RECT 5.680000  8.560000 5.940000  8.630000 ;
        RECT 5.750000  8.630000 6.010000  8.700000 ;
        RECT 5.820000  8.700000 6.080000  8.770000 ;
        RECT 5.890000  8.770000 6.150000  8.840000 ;
        RECT 5.960000  8.840000 6.220000  8.910000 ;
        RECT 5.965000 42.985000 6.225000 43.625000 ;
        RECT 5.970000 42.980000 6.220000 42.985000 ;
        RECT 5.975000 39.420000 6.255000 39.470000 ;
        RECT 5.975000 39.470000 6.205000 39.520000 ;
        RECT 5.975000 39.520000 6.205000 42.965000 ;
        RECT 5.975000 42.965000 6.205000 42.970000 ;
        RECT 5.975000 42.970000 6.210000 42.975000 ;
        RECT 5.975000 42.975000 6.215000 42.980000 ;
        RECT 5.985000 39.410000 6.305000 39.420000 ;
        RECT 6.030000  8.910000 6.290000  8.980000 ;
        RECT 6.055000 39.340000 6.315000 39.410000 ;
        RECT 6.100000  8.980000 6.360000  9.050000 ;
        RECT 6.125000 39.270000 6.385000 39.340000 ;
        RECT 6.170000  9.050000 6.430000  9.120000 ;
        RECT 6.195000 39.200000 6.455000 39.270000 ;
        RECT 6.240000  9.120000 6.500000  9.190000 ;
        RECT 6.265000 39.130000 6.525000 39.200000 ;
        RECT 6.310000  9.190000 6.570000  9.260000 ;
        RECT 6.335000 39.060000 6.595000 39.130000 ;
        RECT 6.380000  9.260000 6.640000  9.330000 ;
        RECT 6.405000 38.990000 6.665000 39.060000 ;
        RECT 6.450000  9.330000 6.710000  9.400000 ;
        RECT 6.475000  9.400000 6.780000  9.425000 ;
        RECT 6.475000 38.920000 6.735000 38.990000 ;
        RECT 6.525000  9.425000 6.805000  9.475000 ;
        RECT 6.525000 38.870000 6.805000 38.920000 ;
        RECT 6.575000  9.475000 6.805000  9.525000 ;
        RECT 6.575000  9.525000 6.805000 38.820000 ;
        RECT 6.575000 38.820000 6.805000 38.870000 ;
    END
  END OE_N
  PIN OUT
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355000  0.000000 22.615000  6.315000 ;
        RECT 22.355000  6.315000 22.615000  6.370000 ;
        RECT 22.355000  6.370000 22.670000  6.425000 ;
        RECT 22.425000  6.425000 22.725000  6.495000 ;
        RECT 22.495000  6.495000 22.795000  6.565000 ;
        RECT 22.565000  6.565000 22.865000  6.635000 ;
        RECT 22.635000  6.635000 22.935000  6.705000 ;
        RECT 22.655000  6.705000 23.005000  6.725000 ;
        RECT 22.710000  6.725000 23.025000  6.780000 ;
        RECT 22.765000  6.780000 23.025000  6.835000 ;
        RECT 22.765000  6.835000 23.025000 14.375000 ;
        RECT 22.765000 14.375000 23.025000 14.430000 ;
        RECT 22.765000 14.430000 23.080000 14.485000 ;
        RECT 22.835000 14.485000 23.135000 14.555000 ;
        RECT 22.905000 14.555000 23.205000 14.625000 ;
        RECT 22.975000 14.625000 23.275000 14.695000 ;
        RECT 23.045000 14.695000 23.345000 14.765000 ;
        RECT 23.095000 38.695000 23.735000 38.955000 ;
        RECT 23.115000 14.765000 23.415000 14.835000 ;
        RECT 23.185000 14.835000 23.485000 14.905000 ;
        RECT 23.255000 14.905000 23.555000 14.975000 ;
        RECT 23.265000 38.625000 23.735000 38.695000 ;
        RECT 23.325000 14.975000 23.625000 15.045000 ;
        RECT 23.335000 38.555000 23.735000 38.625000 ;
        RECT 23.395000 15.045000 23.695000 15.115000 ;
        RECT 23.405000 38.485000 23.735000 38.555000 ;
        RECT 23.465000 15.115000 23.765000 15.185000 ;
        RECT 23.475000 25.180000 23.790000 25.235000 ;
        RECT 23.475000 25.235000 23.735000 25.290000 ;
        RECT 23.475000 25.290000 23.735000 38.415000 ;
        RECT 23.475000 38.415000 23.735000 38.485000 ;
        RECT 23.510000 25.145000 23.845000 25.180000 ;
        RECT 23.535000 15.185000 23.835000 15.255000 ;
        RECT 23.545000 15.255000 23.905000 15.265000 ;
        RECT 23.545000 25.110000 23.880000 25.145000 ;
        RECT 23.600000 15.265000 23.915000 15.320000 ;
        RECT 23.600000 25.055000 23.915000 25.110000 ;
        RECT 23.655000 15.320000 23.915000 15.375000 ;
        RECT 23.655000 15.375000 23.915000 25.000000 ;
        RECT 23.655000 25.000000 23.915000 25.055000 ;
    END
  END OUT
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  216.1550 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.115000 125.470000 53.655000 147.015000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    ANTENNAPARTIALMETALSIDEAREA  3.812250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280000 0.000000 76.920000 1.625000 ;
        RECT 76.280000 1.625000 76.920000 1.695000 ;
        RECT 76.280000 1.695000 76.990000 1.765000 ;
        RECT 76.280000 1.765000 77.060000 1.835000 ;
        RECT 76.280000 1.835000 77.130000 1.905000 ;
        RECT 76.280000 1.905000 77.200000 1.975000 ;
        RECT 76.280000 1.975000 77.270000 2.045000 ;
        RECT 76.280000 2.045000 77.340000 2.055000 ;
        RECT 76.350000 2.055000 77.350000 2.125000 ;
        RECT 76.420000 2.125000 77.420000 2.195000 ;
        RECT 76.490000 2.195000 77.490000 2.265000 ;
        RECT 76.560000 2.265000 77.560000 2.335000 ;
        RECT 76.630000 2.335000 77.630000 2.405000 ;
        RECT 76.700000 2.405000 77.700000 2.475000 ;
        RECT 76.770000 2.475000 77.770000 2.545000 ;
        RECT 76.820000 2.545000 77.840000 2.595000 ;
        RECT 76.890000 2.595000 77.890000 2.665000 ;
        RECT 76.960000 2.665000 77.890000 2.735000 ;
        RECT 77.030000 2.735000 77.890000 2.805000 ;
        RECT 77.100000 2.805000 77.890000 2.875000 ;
        RECT 77.150000 2.875000 77.890000 2.925000 ;
        RECT 77.150000 2.925000 77.890000 5.235000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    ANTENNAPARTIALMETALSIDEAREA  2.618000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275000 0.000000 68.925000 3.960000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    ANTENNAPARTIALCUTAREA  4.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.600000  7.425000 60.560000   7.575000 ;
        RECT 59.600000  7.575000 60.410000   7.725000 ;
        RECT 59.600000  7.725000 60.385000   7.750000 ;
        RECT 59.600000  7.750000 60.385000  10.610000 ;
        RECT 59.600000 10.610000 60.385000  10.760000 ;
        RECT 59.600000 10.760000 60.535000  10.910000 ;
        RECT 59.600000 10.910000 60.685000  10.935000 ;
        RECT 59.655000  7.370000 60.710000   7.425000 ;
        RECT 59.750000 10.935000 60.710000  11.085000 ;
        RECT 59.805000  7.220000 60.765000   7.370000 ;
        RECT 59.900000 11.085000 60.860000  11.235000 ;
        RECT 59.955000  7.070000 60.915000   7.220000 ;
        RECT 59.985000  7.040000 63.890000   7.070000 ;
        RECT 60.050000 11.235000 61.010000  11.385000 ;
        RECT 60.135000  6.890000 63.890000   7.040000 ;
        RECT 60.200000 11.385000 61.160000  11.535000 ;
        RECT 60.285000  6.740000 63.890000   6.890000 ;
        RECT 60.350000 11.535000 61.310000  11.685000 ;
        RECT 60.435000  6.590000 63.890000   6.740000 ;
        RECT 60.500000 11.685000 61.460000  11.835000 ;
        RECT 60.585000  6.440000 63.890000   6.590000 ;
        RECT 60.610000 19.065000 61.570000  19.215000 ;
        RECT 60.610000 19.215000 61.420000  19.365000 ;
        RECT 60.610000 19.365000 61.395000  19.390000 ;
        RECT 60.610000 19.390000 61.395000  47.360000 ;
        RECT 60.650000 11.835000 61.610000  11.985000 ;
        RECT 60.690000 18.985000 61.720000  19.065000 ;
        RECT 60.735000  6.290000 63.890000   6.440000 ;
        RECT 60.800000 11.985000 61.760000  12.135000 ;
        RECT 60.840000 18.835000 61.800000  18.985000 ;
        RECT 60.950000 12.135000 61.910000  12.285000 ;
        RECT 60.990000 18.685000 61.950000  18.835000 ;
        RECT 61.100000 12.285000 62.060000  12.435000 ;
        RECT 61.140000 12.435000 62.210000  12.475000 ;
        RECT 61.140000 18.535000 62.100000  18.685000 ;
        RECT 61.170000 18.505000 62.250000  18.535000 ;
        RECT 61.290000 12.475000 62.250000  12.625000 ;
        RECT 61.320000 18.355000 62.250000  18.505000 ;
        RECT 61.440000 12.625000 62.250000  12.775000 ;
        RECT 61.470000 12.775000 62.250000  12.805000 ;
        RECT 61.470000 12.805000 62.250000  18.205000 ;
        RECT 61.470000 18.205000 62.250000  18.355000 ;
        RECT 61.710000 35.760000 63.070000  35.910000 ;
        RECT 61.710000 35.910000 62.920000  36.060000 ;
        RECT 61.710000 36.060000 62.780000  36.200000 ;
        RECT 61.710000 36.200000 62.780000  73.005000 ;
        RECT 61.710000 73.005000 62.780000  73.155000 ;
        RECT 61.710000 73.155000 62.930000  73.305000 ;
        RECT 61.710000 73.305000 63.080000  73.455000 ;
        RECT 61.710000 73.455000 63.230000  73.605000 ;
        RECT 61.710000 73.605000 63.380000  73.755000 ;
        RECT 61.710000 73.755000 63.530000  73.905000 ;
        RECT 61.710000 73.905000 63.680000  74.055000 ;
        RECT 61.710000 74.055000 63.830000  74.185000 ;
        RECT 61.735000 35.735000 63.220000  35.760000 ;
        RECT 61.750000 74.185000 63.960000  74.225000 ;
        RECT 61.790000 74.225000 64.000000  74.265000 ;
        RECT 61.885000 35.585000 63.245000  35.735000 ;
        RECT 61.940000 74.265000 68.555000  74.415000 ;
        RECT 62.035000 35.435000 63.395000  35.585000 ;
        RECT 62.090000 74.415000 68.705000  74.565000 ;
        RECT 62.185000 35.285000 63.545000  35.435000 ;
        RECT 62.220000  6.155000 63.890000   6.290000 ;
        RECT 62.235000  7.070000 63.890000   7.220000 ;
        RECT 62.240000 74.565000 68.855000  74.715000 ;
        RECT 62.325000 35.145000 63.695000  35.285000 ;
        RECT 62.370000  6.005000 63.890000   6.155000 ;
        RECT 62.385000  7.220000 63.890000   7.370000 ;
        RECT 62.390000 74.715000 69.005000  74.865000 ;
        RECT 62.475000 34.995000 63.695000  35.145000 ;
        RECT 62.520000  5.855000 63.890000   6.005000 ;
        RECT 62.535000  7.370000 63.890000   7.520000 ;
        RECT 62.540000 74.865000 69.155000  75.015000 ;
        RECT 62.625000 17.825000 63.890000  18.070000 ;
        RECT 62.625000 18.070000 63.795000  18.165000 ;
        RECT 62.625000 18.165000 63.700000  18.260000 ;
        RECT 62.625000 18.260000 63.695000  18.265000 ;
        RECT 62.625000 18.265000 63.695000  34.845000 ;
        RECT 62.625000 34.845000 63.695000  34.995000 ;
        RECT 62.630000 17.820000 63.890000  17.825000 ;
        RECT 62.670000  5.705000 63.890000   5.855000 ;
        RECT 62.685000  7.520000 63.890000   7.670000 ;
        RECT 62.690000 75.015000 69.305000  75.165000 ;
        RECT 62.725000 17.725000 63.890000  17.820000 ;
        RECT 62.820000  0.000000 63.890000   5.555000 ;
        RECT 62.820000  5.555000 63.890000   5.705000 ;
        RECT 62.820000  7.670000 63.890000   7.805000 ;
        RECT 62.820000  7.805000 63.890000  17.630000 ;
        RECT 62.820000 17.630000 63.890000  17.725000 ;
        RECT 62.840000 75.165000 69.455000  75.315000 ;
        RECT 62.860000 75.315000 69.605000  75.335000 ;
        RECT 67.870000 75.335000 69.625000  75.400000 ;
        RECT 67.935000 75.400000 69.690000  75.465000 ;
        RECT 67.940000 75.465000 69.755000  75.470000 ;
        RECT 68.090000 75.470000 69.760000  75.620000 ;
        RECT 68.240000 75.620000 69.760000  75.770000 ;
        RECT 68.390000 75.770000 69.760000  75.920000 ;
        RECT 68.540000 75.920000 69.760000  76.070000 ;
        RECT 68.690000 76.070000 69.760000  76.220000 ;
        RECT 68.690000 76.220000 69.760000 101.910000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.000000 106.585000 12.500000 118.955000 ;
        RECT 7.665000 118.955000 12.500000 119.105000 ;
        RECT 7.815000 119.105000 12.500000 119.255000 ;
        RECT 7.850000 106.565000 12.500000 106.585000 ;
        RECT 7.965000 119.255000 12.500000 119.405000 ;
        RECT 8.000000 106.415000 12.500000 106.565000 ;
        RECT 8.115000 119.405000 12.500000 119.555000 ;
        RECT 8.150000 106.265000 12.500000 106.415000 ;
        RECT 8.265000 119.555000 12.500000 119.705000 ;
        RECT 8.300000 106.115000 12.500000 106.265000 ;
        RECT 8.415000 119.705000 12.500000 119.855000 ;
        RECT 8.450000 105.965000 12.500000 106.115000 ;
        RECT 8.565000 119.855000 12.500000 120.005000 ;
        RECT 8.600000 105.815000 12.500000 105.965000 ;
        RECT 8.715000 120.005000 12.500000 120.155000 ;
        RECT 8.750000 105.665000 12.500000 105.815000 ;
        RECT 8.865000 120.155000 12.500000 120.305000 ;
        RECT 8.900000 105.515000 12.500000 105.665000 ;
        RECT 9.015000 120.305000 12.500000 120.455000 ;
        RECT 9.050000 105.365000 12.500000 105.515000 ;
        RECT 9.165000 120.455000 12.500000 120.605000 ;
        RECT 9.200000 105.215000 12.500000 105.365000 ;
        RECT 9.315000 120.605000 12.500000 120.755000 ;
        RECT 9.350000 105.065000 12.500000 105.215000 ;
        RECT 9.465000 120.755000 12.500000 120.905000 ;
        RECT 9.500000 104.915000 12.500000 105.065000 ;
        RECT 9.615000 120.905000 12.500000 121.055000 ;
        RECT 9.650000 104.765000 12.500000 104.915000 ;
        RECT 9.765000 121.055000 12.500000 121.205000 ;
        RECT 9.800000 104.615000 12.500000 104.765000 ;
        RECT 9.810000 121.205000 12.500000 121.250000 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.390000 1.185000 78.210000 1.465000 ;
        RECT 77.470000 1.125000 78.120000 1.185000 ;
        RECT 77.540000 1.055000 78.050000 1.125000 ;
        RECT 77.610000 0.000000 77.870000 0.875000 ;
        RECT 77.610000 0.875000 77.870000 0.930000 ;
        RECT 77.610000 0.930000 77.925000 0.985000 ;
        RECT 77.610000 0.985000 77.980000 1.055000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    ANTENNAPARTIALMETALSIDEAREA  85.19250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.230000 50.760000 76.475000 50.805000 ;
        RECT 76.230000 50.805000 76.430000 50.850000 ;
        RECT 76.230000 50.850000 76.430000 52.425000 ;
        RECT 76.230000 52.425000 76.430000 52.470000 ;
        RECT 76.230000 52.470000 76.475000 52.515000 ;
        RECT 76.280000 50.710000 76.520000 50.760000 ;
        RECT 76.300000 52.515000 76.520000 52.585000 ;
        RECT 76.350000 50.640000 76.570000 50.710000 ;
        RECT 76.370000 52.585000 76.590000 52.655000 ;
        RECT 76.420000 50.570000 76.640000 50.640000 ;
        RECT 76.440000 52.655000 76.660000 52.725000 ;
        RECT 76.490000 50.500000 76.710000 50.570000 ;
        RECT 76.510000 52.725000 76.730000 52.795000 ;
        RECT 76.560000 50.430000 76.780000 50.500000 ;
        RECT 76.580000 52.795000 76.800000 52.865000 ;
        RECT 76.630000 50.360000 76.850000 50.430000 ;
        RECT 76.650000 52.865000 76.870000 52.935000 ;
        RECT 76.700000 50.290000 76.920000 50.360000 ;
        RECT 76.720000 52.935000 76.940000 53.005000 ;
        RECT 76.770000 50.220000 76.990000 50.290000 ;
        RECT 76.790000 53.005000 77.010000 53.075000 ;
        RECT 76.825000 53.075000 77.080000 53.110000 ;
        RECT 76.840000 50.150000 77.060000 50.220000 ;
        RECT 76.870000 53.110000 77.115000 53.155000 ;
        RECT 76.900000 96.210000 77.130000 96.225000 ;
        RECT 76.910000 50.080000 77.130000 50.150000 ;
        RECT 76.915000 53.155000 77.115000 53.200000 ;
        RECT 76.915000 53.200000 77.115000 96.195000 ;
        RECT 76.915000 96.195000 77.115000 96.210000 ;
        RECT 76.980000 50.010000 77.200000 50.080000 ;
        RECT 77.050000 49.940000 77.270000 50.010000 ;
        RECT 77.120000 49.870000 77.340000 49.940000 ;
        RECT 77.190000 49.800000 77.410000 49.870000 ;
        RECT 77.260000 49.730000 77.480000 49.800000 ;
        RECT 77.330000 49.660000 77.550000 49.730000 ;
        RECT 77.400000 49.590000 77.620000 49.660000 ;
        RECT 77.470000 49.520000 77.690000 49.590000 ;
        RECT 77.540000 49.450000 77.760000 49.520000 ;
        RECT 77.610000 49.380000 77.830000 49.450000 ;
        RECT 77.680000 49.310000 77.900000 49.380000 ;
        RECT 77.750000 49.240000 77.970000 49.310000 ;
        RECT 77.820000 49.170000 78.040000 49.240000 ;
        RECT 77.890000 49.100000 78.110000 49.170000 ;
        RECT 77.960000 49.030000 78.180000 49.100000 ;
        RECT 78.030000 48.960000 78.250000 49.030000 ;
        RECT 78.100000 48.890000 78.320000 48.960000 ;
        RECT 78.170000 48.820000 78.390000 48.890000 ;
        RECT 78.240000 48.750000 78.460000 48.820000 ;
        RECT 78.310000 48.680000 78.530000 48.750000 ;
        RECT 78.380000 48.610000 78.600000 48.680000 ;
        RECT 78.450000 48.540000 78.670000 48.610000 ;
        RECT 78.520000 48.470000 78.740000 48.540000 ;
        RECT 78.590000 48.400000 78.810000 48.470000 ;
        RECT 78.615000 10.265000 78.910000 10.340000 ;
        RECT 78.615000 10.340000 78.860000 10.390000 ;
        RECT 78.615000 10.390000 78.810000 10.440000 ;
        RECT 78.615000 10.440000 78.805000 10.445000 ;
        RECT 78.615000 10.445000 78.805000 16.245000 ;
        RECT 78.615000 16.245000 78.805000 16.285000 ;
        RECT 78.615000 16.285000 78.845000 16.325000 ;
        RECT 78.620000 10.260000 78.910000 10.265000 ;
        RECT 78.660000 48.330000 78.880000 48.400000 ;
        RECT 78.665000 10.215000 78.910000 10.260000 ;
        RECT 78.685000 16.325000 78.885000 16.395000 ;
        RECT 78.705000  0.000000 78.905000  1.125000 ;
        RECT 78.705000  1.125000 78.905000  1.130000 ;
        RECT 78.705000  1.130000 78.910000  1.215000 ;
        RECT 78.710000  1.215000 78.910000  1.220000 ;
        RECT 78.710000  1.220000 78.910000 10.170000 ;
        RECT 78.710000 10.170000 78.910000 10.215000 ;
        RECT 78.730000 48.260000 78.950000 48.330000 ;
        RECT 78.755000 16.395000 78.955000 16.465000 ;
        RECT 78.800000 48.190000 79.020000 48.260000 ;
        RECT 78.825000 16.465000 79.025000 16.535000 ;
        RECT 78.870000 48.120000 79.090000 48.190000 ;
        RECT 78.895000 16.535000 79.095000 16.605000 ;
        RECT 78.940000 48.050000 79.160000 48.120000 ;
        RECT 78.965000 16.605000 79.165000 16.675000 ;
        RECT 79.010000 47.980000 79.230000 48.050000 ;
        RECT 79.035000 16.675000 79.235000 16.745000 ;
        RECT 79.080000 47.910000 79.300000 47.980000 ;
        RECT 79.105000 16.745000 79.305000 16.815000 ;
        RECT 79.150000 47.840000 79.370000 47.910000 ;
        RECT 79.175000 16.815000 79.375000 16.885000 ;
        RECT 79.220000 47.770000 79.440000 47.840000 ;
        RECT 79.240000 16.885000 79.445000 16.950000 ;
        RECT 79.270000 47.720000 79.510000 47.770000 ;
        RECT 79.280000 16.950000 79.510000 16.990000 ;
        RECT 79.320000 16.990000 79.510000 17.030000 ;
        RECT 79.320000 17.030000 79.510000 47.670000 ;
        RECT 79.320000 47.670000 79.510000 47.720000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALMETALSIDEAREA  165.2660 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715000 0.000000 79.915000 96.000000 ;
    END
  END TIE_LO_ESD
  PIN VTRIP_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130000 0.000000 6.390000 1.440000 ;
        RECT 6.130000 1.440000 6.390000 1.495000 ;
        RECT 6.130000 1.495000 6.445000 1.550000 ;
        RECT 6.200000 1.550000 6.500000 1.620000 ;
        RECT 6.270000 1.620000 6.570000 1.690000 ;
        RECT 6.340000 1.690000 6.640000 1.760000 ;
        RECT 6.410000 1.760000 6.710000 1.830000 ;
        RECT 6.480000 1.830000 6.780000 1.900000 ;
        RECT 6.550000 1.900000 6.850000 1.970000 ;
        RECT 6.620000 1.970000 6.920000 2.040000 ;
        RECT 6.690000 2.040000 6.990000 2.110000 ;
        RECT 6.760000 2.110000 7.060000 2.180000 ;
        RECT 6.830000 2.180000 7.130000 2.250000 ;
        RECT 6.900000 2.250000 7.200000 2.320000 ;
        RECT 6.970000 2.320000 7.270000 2.390000 ;
        RECT 7.040000 2.390000 7.340000 2.460000 ;
        RECT 7.110000 2.460000 7.410000 2.530000 ;
        RECT 7.180000 2.530000 7.480000 2.600000 ;
        RECT 7.250000 2.600000 7.550000 2.670000 ;
        RECT 7.320000 2.670000 7.620000 2.740000 ;
        RECT 7.390000 2.740000 7.690000 2.810000 ;
        RECT 7.460000 2.810000 7.760000 2.880000 ;
        RECT 7.530000 2.880000 7.830000 2.950000 ;
        RECT 7.600000 2.950000 7.900000 3.020000 ;
        RECT 7.670000 3.020000 7.970000 3.090000 ;
        RECT 7.740000 3.090000 8.040000 3.160000 ;
        RECT 7.810000 3.160000 8.110000 3.230000 ;
        RECT 7.880000 3.230000 8.180000 3.300000 ;
        RECT 7.950000 3.300000 8.250000 3.370000 ;
        RECT 8.020000 3.370000 8.320000 3.440000 ;
        RECT 8.090000 3.440000 8.390000 3.510000 ;
        RECT 8.160000 3.510000 8.460000 3.580000 ;
        RECT 8.230000 3.580000 8.530000 3.650000 ;
        RECT 8.300000 3.650000 8.600000 3.720000 ;
        RECT 8.335000 3.720000 8.670000 3.755000 ;
        RECT 8.390000 3.755000 8.705000 3.810000 ;
        RECT 8.445000 3.810000 8.705000 3.865000 ;
        RECT 8.445000 3.865000 8.705000 6.780000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 8.885000 80.000000 13.535000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 2.035000 80.000000 7.485000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.035000 14.935000 80.000000 18.385000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 19.785000 80.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 70.035000 80.000000 95.000000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 64.085000 80.000000 68.535000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 36.735000 80.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 47.735000 80.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 51.645000 80.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 56.405000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 41.585000 80.000000 46.235000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 175.785000 80.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 25.835000 80.000000 30.485000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 58.235000 80.000000 62.685000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 31.885000 80.000000 35.335000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.115000  95.895000 45.710000  95.955000 ;
      RECT -0.115000  95.955000  4.915000 130.220000 ;
      RECT -0.115000 131.275000  4.915000 140.050000 ;
      RECT -0.115000 140.050000  1.495000 140.150000 ;
      RECT -0.115000 145.155000  1.495000 145.210000 ;
      RECT -0.115000 145.210000  4.915000 170.090000 ;
      RECT -0.085000  93.065000  9.000000  95.255000 ;
      RECT -0.085000  95.255000 45.710000  95.895000 ;
      RECT -0.085000 130.220000  4.915000 130.225000 ;
      RECT -0.085000 130.995000  4.915000 131.275000 ;
      RECT -0.085000 170.090000  4.915000 178.645000 ;
      RECT  0.950000  18.885000  1.310000  19.055000 ;
      RECT  0.980000  21.465000  1.310000  21.635000 ;
      RECT  1.120000  22.325000  1.310000  22.495000 ;
      RECT  1.150000  19.745000  1.310000  19.915000 ;
      RECT  1.150000  20.605000  1.310000  20.775000 ;
      RECT  1.690000  45.545000  4.585000  45.715000 ;
      RECT  2.260000 145.155000  4.700000 145.210000 ;
      RECT  5.875000   5.940000  6.405000   6.465000 ;
      RECT  6.490000  88.950000  9.000000  93.065000 ;
      RECT  7.805000   5.400000 67.100000   6.230000 ;
      RECT  9.300000  32.000000  9.660000  36.750000 ;
      RECT 10.330000  32.000000 10.690000  36.750000 ;
      RECT 11.410000  32.000000 11.665000  37.260000 ;
      RECT 11.940000  31.110000 12.365000  36.765000 ;
      RECT 12.610000  32.000000 13.140000  37.260000 ;
      RECT 13.390000  32.000000 13.920000  36.750000 ;
      RECT 14.170000  32.000000 14.700000  36.750000 ;
      RECT 14.170000  36.750000 14.305000  37.260000 ;
      RECT 14.320000  26.760000 14.500000  29.470000 ;
      RECT 14.320000  29.470000 14.670000  29.570000 ;
      RECT 14.320000  29.570000 14.490000  30.110000 ;
      RECT 14.955000  32.000000 15.485000  37.260000 ;
      RECT 15.105000  26.760000 15.635000  29.690000 ;
      RECT 15.730000  32.000000 16.260000  36.750000 ;
      RECT 15.730000 179.435000 68.925000 179.450000 ;
      RECT 15.730000 179.450000 77.885000 179.980000 ;
      RECT 15.730000 179.980000 68.925000 180.205000 ;
      RECT 15.885000  26.760000 16.415000  29.470000 ;
      RECT 16.510000  32.000000 16.950000  37.260000 ;
      RECT 16.670000  26.760000 17.200000  29.690000 ;
      RECT 17.210000  32.000000 17.650000  36.750000 ;
      RECT 18.035000  26.760000 18.450000  29.470000 ;
      RECT 18.140000  32.060000 18.630000  36.750000 ;
      RECT 19.040000  26.760000 19.455000  29.470000 ;
      RECT 19.050000  32.000000 19.580000  36.750000 ;
      RECT 19.790000  26.760000 20.320000  29.470000 ;
      RECT 20.640000  32.000000 21.170000  36.750000 ;
      RECT 21.690000  26.760000 22.130000  29.470000 ;
      RECT 22.170000  32.000000 22.700000  36.755000 ;
      RECT 23.725000  32.000000 24.255000  36.755000 ;
      RECT 23.800000  26.760000 24.160000  29.470000 ;
      RECT 24.340000  25.580000 26.330000  25.905000 ;
      RECT 24.340000  25.905000 24.835000  29.690000 ;
      RECT 25.015000  26.760000 25.545000  29.470000 ;
      RECT 25.675000  32.250000 26.090000  37.000000 ;
      RECT 25.930000  59.095000 28.100000  60.125000 ;
      RECT 25.935000  57.585000 29.370000  58.865000 ;
      RECT 26.225000  19.595000 26.670000  24.375000 ;
      RECT 26.385000  32.250000 26.865000  37.330000 ;
      RECT 26.390000  26.760000 26.750000  29.690000 ;
      RECT 26.525000  67.105000 29.670000  67.815000 ;
      RECT 26.975000  19.600000 27.420000  24.365000 ;
      RECT 27.045000  32.250000 27.575000  37.000000 ;
      RECT 27.490000  63.970000 29.315000  64.550000 ;
      RECT 27.510000  26.490000 28.090000  30.360000 ;
      RECT 27.675000  68.735000 29.670000  69.445000 ;
      RECT 27.830000  32.245000 28.360000  37.330000 ;
      RECT 28.340000  59.180000 28.510000  59.710000 ;
      RECT 28.605000  32.250000 29.135000  37.005000 ;
      RECT 28.680000  18.995000 29.210000  23.750000 ;
      RECT 28.860000  95.125000 45.710000  95.255000 ;
      RECT 29.035000  56.755000 29.565000  57.285000 ;
      RECT 29.390000  18.965000 30.080000  23.745000 ;
      RECT 29.390000  32.250000 29.920000  37.330000 ;
      RECT 30.165000  32.250000 30.695000  37.000000 ;
      RECT 30.270000  18.995000 30.800000  23.745000 ;
      RECT 30.950000  32.250000 31.375000  37.330000 ;
      RECT 31.660000  32.250000 32.085000  37.005000 ;
      RECT 31.820000  18.995000 32.350000  23.745000 ;
      RECT 32.410000  32.060000 33.070000  36.750000 ;
      RECT 33.500000  31.990000 33.930000  37.080000 ;
      RECT 34.305000  31.975000 34.865000  36.750000 ;
      RECT 35.060000  31.990000 35.490000  37.080000 ;
      RECT 35.865000  31.975000 36.425000  36.750000 ;
      RECT 35.870000  26.885000 36.305000  28.235000 ;
      RECT 36.620000  31.990000 37.050000  37.080000 ;
      RECT 37.425000  31.975000 37.985000  36.750000 ;
      RECT 38.180000  31.990000 38.610000  37.080000 ;
      RECT 38.985000  31.975000 39.545000  36.750000 ;
      RECT 39.270000  26.885000 39.690000  28.235000 ;
      RECT 39.685000  95.955000 45.710000  96.105000 ;
      RECT 39.715000  31.990000 40.090000  36.750000 ;
      RECT 40.580000  32.155000 40.900000  36.710000 ;
      RECT 43.380000  24.850000 43.870000  27.560000 ;
      RECT 43.855000 180.205000 44.500000 180.370000 ;
      RECT 44.200000  33.270000 44.390000  36.510000 ;
      RECT 45.310000  36.340000 46.360000  36.970000 ;
      RECT 49.340000  32.065000 51.760000  32.445000 ;
      RECT 51.105000  32.445000 51.760000  33.690000 ;
      RECT 52.050000  24.855000 52.580000  27.565000 ;
      RECT 53.470000  24.855000 54.000000  27.565000 ;
      RECT 54.870000  24.855000 55.400000  27.565000 ;
      RECT 56.725000 180.205000 57.305000 180.370000 ;
      RECT 59.360000   2.260000 59.720000   3.430000 ;
      RECT 61.115000   5.230000 67.290000   5.345000 ;
      RECT 61.115000   5.345000 67.100000   5.400000 ;
      RECT 61.370000   5.080000 67.290000   5.230000 ;
      RECT 61.560000   4.765000 67.290000   5.080000 ;
      RECT 64.375000   0.250000 66.075000   1.000000 ;
      RECT 65.660000   6.230000 67.100000   9.570000 ;
      RECT 66.390000   9.570000 67.100000   9.575000 ;
      RECT 66.390000   9.575000 69.665000   9.745000 ;
      RECT 66.390000   9.745000 71.650000  10.185000 ;
      RECT 68.290000   1.940000 69.255000   3.960000 ;
      RECT 69.165000 128.445000 79.585000 130.115000 ;
      RECT 69.625000 179.435000 77.885000 179.450000 ;
      RECT 69.625000 179.980000 77.885000 180.205000 ;
      RECT 69.665000  10.185000 71.650000  11.425000 ;
      RECT 72.315000   1.940000 74.335000   4.420000 ;
      RECT 73.080000   8.080000 74.910000   8.830000 ;
      RECT 74.910000   5.170000 76.930000   5.800000 ;
      RECT 74.910000   5.800000 79.430000   7.820000 ;
      RECT 77.195000   3.705000 79.430000   4.420000 ;
      RECT 77.195000   4.420000 77.775000   5.170000 ;
      RECT 77.410000   3.700000 79.430000   3.705000 ;
      RECT 77.410000   7.820000 79.430000   8.080000 ;
      RECT 79.880000  19.485000 80.120000  25.015000 ;
      RECT 79.880000  30.115000 80.120000  35.725000 ;
    LAYER met1 ;
      RECT -0.115000  95.895000  1.495000 130.220000 ;
      RECT -0.115000 131.275000  1.495000 170.090000 ;
      RECT  0.000000   0.000000  5.565000   1.560000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000 62.290000   2.055000 ;
      RECT  0.000000   1.560000  5.565000   1.565000 ;
      RECT  0.000000   1.565000  5.565000   2.055000 ;
      RECT  0.000000   1.565000 35.574000   1.635000 ;
      RECT  0.000000   1.635000 35.504000   1.705000 ;
      RECT  0.000000   1.705000 35.434000   1.775000 ;
      RECT  0.000000   1.775000 35.364000   1.845000 ;
      RECT  0.000000   1.845000 35.294000   1.915000 ;
      RECT  0.000000   1.915000 35.224000   1.985000 ;
      RECT  0.000000   1.985000 35.154000   2.055000 ;
      RECT  0.000000   2.055000  5.565000   2.875000 ;
      RECT  0.000000   2.055000 80.000000 106.585000 ;
      RECT  0.000000   2.875000 11.260000   3.155000 ;
      RECT  0.000000   3.155000 67.995000   4.240000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   4.240000 76.885000   5.515000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   5.515000 80.000000  10.335000 ;
      RECT  0.000000  10.335000  1.340000  11.155000 ;
      RECT  0.000000  11.155000  0.750000  12.425000 ;
      RECT  0.000000  12.425000 80.000000  13.120000 ;
      RECT  0.000000  14.320000 76.495000  23.851000 ;
      RECT  0.000000  14.320000 80.000000  16.455000 ;
      RECT  0.000000  17.275000 78.550000  23.851000 ;
      RECT  0.000000  17.275000 78.550000  29.840000 ;
      RECT  0.000000  17.275000 79.605000  19.205000 ;
      RECT  0.000000  17.275000 79.605000  20.649000 ;
      RECT  0.000000  17.275000 79.605000  20.649000 ;
      RECT  0.000000  19.205000 79.605000  20.649000 ;
      RECT  0.000000  20.649000 78.550000  29.840000 ;
      RECT  0.000000  20.649000 79.534000  20.720000 ;
      RECT  0.000000  20.649000 79.534000  20.720000 ;
      RECT  0.000000  20.720000 79.464000  20.790000 ;
      RECT  0.000000  20.720000 79.464000  20.790000 ;
      RECT  0.000000  20.790000 79.394000  20.860000 ;
      RECT  0.000000  20.790000 79.394000  20.860000 ;
      RECT  0.000000  20.860000 79.324000  20.930000 ;
      RECT  0.000000  20.860000 79.324000  20.930000 ;
      RECT  0.000000  20.930000 79.254000  21.000000 ;
      RECT  0.000000  20.930000 79.254000  21.000000 ;
      RECT  0.000000  21.000000 79.184000  21.070000 ;
      RECT  0.000000  21.000000 79.184000  21.070000 ;
      RECT  0.000000  21.070000 79.159000  21.095000 ;
      RECT  0.000000  21.070000 79.159000  21.095000 ;
      RECT  0.000000  23.405000 79.159000  23.475000 ;
      RECT  0.000000  23.405000 79.159000  23.475000 ;
      RECT  0.000000  23.475000 79.229000  23.545000 ;
      RECT  0.000000  23.475000 79.229000  23.545000 ;
      RECT  0.000000  23.545000 79.299000  23.615000 ;
      RECT  0.000000  23.545000 79.299000  23.615000 ;
      RECT  0.000000  23.615000 79.369000  23.685000 ;
      RECT  0.000000  23.615000 79.369000  23.685000 ;
      RECT  0.000000  23.685000 79.439000  23.755000 ;
      RECT  0.000000  23.685000 79.439000  23.755000 ;
      RECT  0.000000  23.755000 79.509000  23.825000 ;
      RECT  0.000000  23.755000 79.509000  23.825000 ;
      RECT  0.000000  23.825000 79.579000  23.850000 ;
      RECT  0.000000  23.825000 79.579000  23.850000 ;
      RECT  0.000000  23.851000 79.605000  25.295000 ;
      RECT  0.000000  25.295000 78.845000  36.005000 ;
      RECT  0.000000  25.295000 78.845000  42.035000 ;
      RECT  0.000000  25.295000 80.000000  29.840000 ;
      RECT  0.000000  29.840000 78.845000  42.035000 ;
      RECT  0.000000  29.840000 79.605000  31.399000 ;
      RECT  0.000000  31.399000 79.534000  31.470000 ;
      RECT  0.000000  31.399000 79.534000  31.470000 ;
      RECT  0.000000  31.470000 79.464000  31.540000 ;
      RECT  0.000000  31.470000 79.464000  31.540000 ;
      RECT  0.000000  31.540000 79.394000  31.610000 ;
      RECT  0.000000  31.540000 79.394000  31.610000 ;
      RECT  0.000000  31.610000 79.324000  31.680000 ;
      RECT  0.000000  31.610000 79.324000  31.680000 ;
      RECT  0.000000  31.680000 79.279000  31.725000 ;
      RECT  0.000000  31.680000 79.279000  31.725000 ;
      RECT  0.000000  31.725000 78.845000  34.115000 ;
      RECT  0.000000  34.115000 79.279000  34.185000 ;
      RECT  0.000000  34.115000 79.279000  34.185000 ;
      RECT  0.000000  34.185000 79.349000  34.255000 ;
      RECT  0.000000  34.185000 79.349000  34.255000 ;
      RECT  0.000000  34.255000 79.419000  34.325000 ;
      RECT  0.000000  34.255000 79.419000  34.325000 ;
      RECT  0.000000  34.325000 79.489000  34.395000 ;
      RECT  0.000000  34.325000 79.489000  34.395000 ;
      RECT  0.000000  34.395000 79.559000  34.440000 ;
      RECT  0.000000  34.395000 79.559000  34.440000 ;
      RECT  0.000000  34.441000 79.605000  36.005000 ;
      RECT  0.000000  36.005000 80.000000  42.035000 ;
      RECT  0.000000  42.035000 78.635000  42.339000 ;
      RECT  0.000000  42.339000 78.564000  42.410000 ;
      RECT  0.000000  42.339000 78.564000  42.410000 ;
      RECT  0.000000  42.410000 78.494000  42.480000 ;
      RECT  0.000000  42.410000 78.494000  42.480000 ;
      RECT  0.000000  42.480000 78.424000  42.550000 ;
      RECT  0.000000  42.480000 78.424000  42.550000 ;
      RECT  0.000000  42.550000 78.354000  42.620000 ;
      RECT  0.000000  42.550000 78.354000  42.620000 ;
      RECT  0.000000  42.620000 78.284000  42.690000 ;
      RECT  0.000000  42.620000 78.284000  42.690000 ;
      RECT  0.000000  42.690000 78.214000  42.760000 ;
      RECT  0.000000  42.690000 78.214000  42.760000 ;
      RECT  0.000000  42.760000 78.144000  42.830000 ;
      RECT  0.000000  42.760000 78.144000  42.830000 ;
      RECT  0.000000  42.830000 78.074000  42.900000 ;
      RECT  0.000000  42.830000 78.074000  42.900000 ;
      RECT  0.000000  42.900000 78.004000  42.970000 ;
      RECT  0.000000  42.900000 78.004000  42.970000 ;
      RECT  0.000000  42.970000 77.999000  42.975000 ;
      RECT  0.000000  42.970000 77.999000  42.975000 ;
      RECT  0.000000  42.975000 78.635000  43.235000 ;
      RECT  0.000000  43.235000 80.000000  44.355000 ;
      RECT  0.000000  44.355000  1.020000  45.010000 ;
      RECT  0.000000  45.010000  0.965000  45.239000 ;
      RECT  0.000000  45.239000  0.894000  45.310000 ;
      RECT  0.000000  45.310000  0.824000  45.380000 ;
      RECT  0.000000  45.380000  0.754000  45.450000 ;
      RECT  0.000000  45.450000  0.684000  45.520000 ;
      RECT  0.000000  45.520000  0.614000  45.590000 ;
      RECT  0.000000  45.590000  0.544000  45.660000 ;
      RECT  0.000000  45.660000  0.474000  45.730000 ;
      RECT  0.000000  45.730000  0.404000  45.800000 ;
      RECT  0.000000  45.800000  0.334000  45.870000 ;
      RECT  0.000000  45.870000  0.264000  45.940000 ;
      RECT  0.000000  45.940000  0.194000  46.010000 ;
      RECT  0.000000  46.010000  0.124000  46.080000 ;
      RECT  0.000000  46.080000  0.054000  46.150000 ;
      RECT  0.000000  46.445000  0.965000  46.580000 ;
      RECT  0.000000  46.580000  1.050000  47.350000 ;
      RECT  0.000000  47.350000 80.000000  93.020000 ;
      RECT  0.000000  93.020000  1.070000  94.660000 ;
      RECT  0.000000  94.660000 11.550000  94.830000 ;
      RECT  0.000000  94.830000  1.985000  95.615000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 130.500000  4.530000 130.715000 ;
      RECT  0.000000 130.715000  1.980000 130.995000 ;
      RECT  0.000000 170.370000  1.980000 178.680000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 80.000000 179.140000 ;
      RECT  0.000000 179.140000 15.445000 180.290000 ;
      RECT  0.000000 180.290000 15.490000 200.000000 ;
      RECT  0.000000 180.290000 80.000000 198.405000 ;
      RECT  0.000000 198.405000 15.490000 200.000000 ;
      RECT  0.210000  13.400000  0.470000  14.040000 ;
      RECT  0.475000  46.125000  5.000000  46.165000 ;
      RECT  0.545000  46.055000  5.000000  46.125000 ;
      RECT  0.615000  45.985000  5.000000  46.055000 ;
      RECT  0.685000  45.915000  5.000000  45.985000 ;
      RECT  0.750000  11.155000 76.825000  12.425000 ;
      RECT  0.750000  13.120000 80.000000  16.125000 ;
      RECT  0.755000  45.845000  5.000000  45.915000 ;
      RECT  0.825000  45.775000  5.000000  45.845000 ;
      RECT  0.895000  45.705000  5.000000  45.775000 ;
      RECT  0.965000  45.635000  5.000000  45.705000 ;
      RECT  1.035000  45.565000  5.000000  45.635000 ;
      RECT  1.105000  45.495000  5.000000  45.565000 ;
      RECT  1.175000  45.425000  5.000000  45.495000 ;
      RECT  1.245000  45.290000  5.000000  45.355000 ;
      RECT  1.245000  45.355000  5.000000  45.425000 ;
      RECT  1.245000  46.165000  5.000000  46.300000 ;
      RECT  1.300000  44.635000  1.730000  45.290000 ;
      RECT  1.330000  46.300000  2.790000  47.070000 ;
      RECT  1.350000  93.300000  8.265000  94.380000 ;
      RECT  1.620000  10.615000  4.025000  10.875000 ;
      RECT  1.775000  95.615000  1.985000 106.585000 ;
      RECT  1.775000 118.955000  1.985000 130.500000 ;
      RECT  1.775000 130.995000  1.980000 140.430000 ;
      RECT  1.775000 140.430000 80.000000 144.875000 ;
      RECT  1.775000 144.875000  1.980000 170.370000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  2.010000  44.355000 80.000000  45.010000 ;
      RECT  2.260000 130.995000  4.700000 139.510000 ;
      RECT  2.260000 139.510000  4.855000 140.150000 ;
      RECT  2.260000 145.155000  4.700000 178.400000 ;
      RECT  2.265000  95.110000  8.970000  95.900000 ;
      RECT  2.265000  95.900000  4.250000 130.220000 ;
      RECT  3.070000  46.580000 80.000000  47.350000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  4.305000   8.145000 80.000000  11.150000 ;
      RECT  4.305000  11.150000 76.825000  11.155000 ;
      RECT  4.530000  96.180000 80.000000 127.980000 ;
      RECT  4.530000 125.130000 70.100000 128.135000 ;
      RECT  4.530000 128.135000 68.825000 130.425000 ;
      RECT  4.530000 130.425000 70.100000 130.500000 ;
      RECT  4.530000 130.500000 80.000000 130.715000 ;
      RECT  4.980000 130.715000 80.000000 139.230000 ;
      RECT  4.980000 144.875000 80.000000 178.680000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  5.135000 139.230000 80.000000 140.430000 ;
      RECT  5.135000 139.230000 80.000000 144.875000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  47.350000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  45.010000 80.000000  46.580000 ;
      RECT  5.565000   0.000000  6.890000   1.560000 ;
      RECT  5.565000   1.560000 22.990000   1.565000 ;
      RECT  5.845000   2.335000 10.120000   2.595000 ;
      RECT  7.170000   0.270000 10.715000   1.280000 ;
      RECT  8.545000  93.020000 11.550000  94.660000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT 10.400000   2.055000 35.084000   2.125000 ;
      RECT 10.400000   2.125000 35.014000   2.195000 ;
      RECT 10.400000   2.195000 34.944000   2.265000 ;
      RECT 10.400000   2.265000 34.879000   2.330000 ;
      RECT 10.400000   2.330000 13.639000   2.335000 ;
      RECT 10.400000   2.335000 11.260000   2.875000 ;
      RECT 10.995000   0.000000 18.955000   1.560000 ;
      RECT 11.540000   2.615000 35.170000   2.685000 ;
      RECT 11.540000   2.685000 35.100000   2.755000 ;
      RECT 11.540000   2.755000 35.070000   2.785000 ;
      RECT 11.540000   2.785000 18.385000   2.790000 ;
      RECT 11.540000   2.790000 13.990000   2.795000 ;
      RECT 11.540000   2.795000 13.985000   2.800000 ;
      RECT 11.540000   2.800000 12.220000   2.835000 ;
      RECT 11.540000   2.835000 12.185000   2.870000 ;
      RECT 11.540000   2.870000 12.180000   2.875000 ;
      RECT 12.301000   3.150000 67.995000   3.155000 ;
      RECT 12.301000   3.150000 67.995000   3.155000 ;
      RECT 12.311000   3.140000 67.995000   3.150000 ;
      RECT 12.311000   3.140000 67.995000   3.150000 ;
      RECT 12.321000   3.130000 67.995000   3.140000 ;
      RECT 12.321000   3.130000 67.995000   3.140000 ;
      RECT 12.346000   3.105000 59.170000   3.130000 ;
      RECT 12.346000   3.105000 59.170000   3.130000 ;
      RECT 12.371000   3.080000 59.170000   3.105000 ;
      RECT 12.371000   3.080000 59.170000   3.105000 ;
      RECT 13.760000   2.610000 35.240000   2.615000 ;
      RECT 14.106000   3.075000 59.170000   3.080000 ;
      RECT 14.106000   3.075000 59.170000   3.080000 ;
      RECT 14.111000   3.070000 59.170000   3.075000 ;
      RECT 14.111000   3.070000 59.170000   3.075000 ;
      RECT 15.725000 179.420000 77.705000 180.010000 ;
      RECT 15.770000 198.685000 56.715000 199.975000 ;
      RECT 18.506000   3.065000 19.369000   3.070000 ;
      RECT 19.235000   0.270000 21.375000   1.280000 ;
      RECT 19.490000   2.785000 28.955000   2.790000 ;
      RECT 21.655000   0.000000 22.990000   1.560000 ;
      RECT 23.270000   0.275000 26.265000   1.285000 ;
      RECT 26.545000   0.000000 33.120000   1.560000 ;
      RECT 26.545000   1.560000 34.265000   1.565000 ;
      RECT 29.076000   3.065000 30.424000   3.070000 ;
      RECT 29.076000   3.065000 30.424000   3.070000 ;
      RECT 30.545000   2.785000 35.065000   2.790000 ;
      RECT 33.400000   0.270000 37.775000   1.280000 ;
      RECT 34.545000   1.280000 37.775000   1.285000 ;
      RECT 35.055000   2.550000 35.245000   2.610000 ;
      RECT 35.125000   2.480000 35.305000   2.550000 ;
      RECT 35.195000   2.410000 35.375000   2.480000 ;
      RECT 35.206000   3.045000 59.170000   3.070000 ;
      RECT 35.206000   3.045000 59.170000   3.070000 ;
      RECT 35.265000   2.340000 35.445000   2.410000 ;
      RECT 35.276000   2.975000 59.170000   3.045000 ;
      RECT 35.276000   2.975000 59.170000   3.045000 ;
      RECT 35.335000   2.270000 35.515000   2.340000 ;
      RECT 35.346000   2.905000 59.170000   2.975000 ;
      RECT 35.346000   2.905000 59.170000   2.975000 ;
      RECT 35.405000   2.200000 35.585000   2.270000 ;
      RECT 35.416000   2.835000 59.170000   2.905000 ;
      RECT 35.416000   2.835000 59.170000   2.905000 ;
      RECT 35.475000   2.130000 35.655000   2.200000 ;
      RECT 35.486000   2.765000 59.170000   2.835000 ;
      RECT 35.486000   2.765000 59.170000   2.835000 ;
      RECT 35.515000   2.090000 43.035000   2.130000 ;
      RECT 35.556000   2.695000 59.170000   2.765000 ;
      RECT 35.556000   2.695000 59.170000   2.765000 ;
      RECT 35.561000   2.690000 42.989000   2.695000 ;
      RECT 35.561000   2.690000 42.989000   2.695000 ;
      RECT 35.585000   2.020000 42.965000   2.090000 ;
      RECT 35.631000   2.620000 42.919000   2.690000 ;
      RECT 35.631000   2.620000 42.919000   2.690000 ;
      RECT 35.655000   1.950000 42.895000   2.020000 ;
      RECT 35.701000   2.550000 42.849000   2.620000 ;
      RECT 35.701000   2.550000 42.849000   2.620000 ;
      RECT 35.771000   2.480000 42.779000   2.550000 ;
      RECT 35.771000   2.480000 42.779000   2.550000 ;
      RECT 35.841000   2.410000 42.709000   2.480000 ;
      RECT 35.841000   2.410000 42.709000   2.480000 ;
      RECT 38.055000   0.000000 40.785000   1.145000 ;
      RECT 38.055000   1.145000 39.110000   1.670000 ;
      RECT 39.390000   1.425000 43.110000   1.495000 ;
      RECT 39.390000   1.495000 43.180000   1.565000 ;
      RECT 39.390000   1.565000 43.250000   1.635000 ;
      RECT 39.390000   1.635000 43.320000   1.685000 ;
      RECT 41.065000   0.270000 41.935000   1.285000 ;
      RECT 42.215000   0.000000 55.320000   1.145000 ;
      RECT 42.875000   2.130000 43.075000   2.180000 ;
      RECT 42.925000   2.180000 43.125000   2.230000 ;
      RECT 42.930000   2.230000 43.175000   2.235000 ;
      RECT 43.000000   2.235000 51.520000   2.305000 ;
      RECT 43.070000   2.305000 51.520000   2.375000 ;
      RECT 43.110000   1.685000 43.370000   1.755000 ;
      RECT 43.110000   2.375000 51.520000   2.415000 ;
      RECT 43.180000   1.755000 43.440000   1.825000 ;
      RECT 43.200000   1.825000 43.510000   1.845000 ;
      RECT 43.270000   1.845000 47.840000   1.915000 ;
      RECT 43.271000   1.145000 62.150000   1.190000 ;
      RECT 43.316000   1.190000 62.150000   1.235000 ;
      RECT 43.340000   1.915000 47.770000   1.985000 ;
      RECT 43.386000   1.235000 47.724000   1.305000 ;
      RECT 43.410000   1.985000 47.700000   2.055000 ;
      RECT 43.430000   2.055000 47.680000   2.075000 ;
      RECT 43.456000   1.305000 47.654000   1.375000 ;
      RECT 43.526000   1.375000 47.584000   1.445000 ;
      RECT 43.596000   1.445000 47.514000   1.515000 ;
      RECT 43.646000   1.515000 47.464000   1.565000 ;
      RECT 47.630000   1.795000 47.910000   1.845000 ;
      RECT 47.680000   1.745000 47.960000   1.795000 ;
      RECT 47.700000   1.725000 55.040000   1.745000 ;
      RECT 47.770000   1.655000 55.040000   1.725000 ;
      RECT 47.840000   1.585000 55.040000   1.655000 ;
      RECT 47.910000   1.515000 55.040000   1.585000 ;
      RECT 50.840000   2.195000 51.520000   2.235000 ;
      RECT 50.880000   2.155000 51.520000   2.195000 ;
      RECT 51.800000   2.025000 54.524000   2.095000 ;
      RECT 51.800000   2.025000 54.524000   2.095000 ;
      RECT 51.800000   2.095000 54.594000   2.165000 ;
      RECT 51.800000   2.095000 54.594000   2.165000 ;
      RECT 51.800000   2.165000 54.664000   2.235000 ;
      RECT 51.800000   2.165000 54.664000   2.235000 ;
      RECT 51.800000   2.235000 54.734000   2.305000 ;
      RECT 51.800000   2.235000 54.734000   2.305000 ;
      RECT 51.800000   2.305000 54.804000   2.375000 ;
      RECT 51.800000   2.305000 54.804000   2.375000 ;
      RECT 51.800000   2.375000 54.874000   2.445000 ;
      RECT 51.800000   2.375000 54.874000   2.445000 ;
      RECT 51.800000   2.445000 54.944000   2.515000 ;
      RECT 51.800000   2.445000 54.944000   2.515000 ;
      RECT 51.800000   2.515000 55.014000   2.585000 ;
      RECT 51.800000   2.515000 55.014000   2.585000 ;
      RECT 51.800000   2.585000 55.084000   2.655000 ;
      RECT 51.800000   2.585000 55.084000   2.655000 ;
      RECT 51.800000   2.656000 59.170000   2.695000 ;
      RECT 54.655000   1.745000 55.040000   1.760000 ;
      RECT 54.670000   1.760000 55.040000   1.775000 ;
      RECT 54.675000   1.775000 55.040000   1.780000 ;
      RECT 54.745000   1.780000 54.875000   1.850000 ;
      RECT 54.815000   1.850000 54.875000   1.920000 ;
      RECT 55.155000   2.060000 59.170000   2.656000 ;
      RECT 55.320000   0.000000 59.170000   1.145000 ;
      RECT 55.320000   1.145000 59.170000   1.235000 ;
      RECT 55.320000   1.235000 59.170000   1.920000 ;
      RECT 55.320000   1.920000 59.170000   2.060000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 198.405000 80.000000 198.420000 ;
      RECT 56.995000 198.420000 71.715000 200.000000 ;
      RECT 59.170000   0.000000 62.150000   1.145000 ;
      RECT 59.170000   1.235000 62.150000   1.920000 ;
      RECT 59.450000   2.200000 59.710000   2.850000 ;
      RECT 59.990000   1.920000 62.150000   2.195000 ;
      RECT 59.990000   2.195000 67.995000   3.130000 ;
      RECT 62.830000   0.000000 80.000000   2.055000 ;
      RECT 62.970000   0.000000 64.095000   1.190000 ;
      RECT 62.970000   1.190000 67.995000   1.960000 ;
      RECT 62.970000   1.960000 67.995000   2.195000 ;
      RECT 64.375000   0.260000 67.295000   0.910000 ;
      RECT 67.575000   0.000000 69.205000   1.190000 ;
      RECT 67.995000   1.190000 69.205000   1.960000 ;
      RECT 68.275000   2.240000 68.925000   3.960000 ;
      RECT 69.105000 128.415000 80.145000 130.145000 ;
      RECT 69.205000   0.000000 80.000000   1.190000 ;
      RECT 69.205000   1.190000 80.000000   1.960000 ;
      RECT 69.205000   1.960000 80.000000   3.365000 ;
      RECT 69.205000   3.365000 76.885000   4.240000 ;
      RECT 70.380000 128.260000 80.145000 128.415000 ;
      RECT 70.380000 130.145000 80.145000 130.220000 ;
      RECT 71.995000 198.700000 76.855000 200.000000 ;
      RECT 76.775000  16.735000 77.415000  16.995000 ;
      RECT 77.105000  11.430000 77.365000  12.145000 ;
      RECT 77.135000 198.420000 80.000000 200.000000 ;
      RECT 77.165000   3.645000 77.805000   5.235000 ;
      RECT 77.645000  11.150000 80.000000  12.425000 ;
      RECT 77.695000  16.455000 80.000000  17.275000 ;
      RECT 77.985000 179.140000 80.000000 180.290000 ;
      RECT 78.085000   3.365000 80.000000   5.515000 ;
      RECT 78.705000  42.665000 79.175000  42.695000 ;
      RECT 78.775000  42.595000 79.175000  42.665000 ;
      RECT 78.830000  21.375000 80.115000  23.125000 ;
      RECT 78.845000  42.525000 79.175000  42.595000 ;
      RECT 78.915000  42.315000 79.175000  42.455000 ;
      RECT 78.915000  42.455000 79.175000  42.525000 ;
      RECT 78.915000  42.695000 79.175000  42.955000 ;
      RECT 79.125000  32.005000 80.115000  33.835000 ;
      RECT 79.325000  21.325000 80.115000  21.375000 ;
      RECT 79.345000  23.125000 80.115000  23.195000 ;
      RECT 79.395000  21.255000 80.115000  21.325000 ;
      RECT 79.415000  23.195000 80.115000  23.265000 ;
      RECT 79.455000  42.035000 80.000000  43.235000 ;
      RECT 79.465000  21.185000 80.115000  21.255000 ;
      RECT 79.465000  31.935000 80.115000  32.005000 ;
      RECT 79.465000  33.835000 80.115000  33.905000 ;
      RECT 79.485000  23.265000 80.115000  23.335000 ;
      RECT 79.535000  21.115000 80.115000  21.185000 ;
      RECT 79.535000  31.865000 80.115000  31.935000 ;
      RECT 79.535000  33.905000 80.115000  33.975000 ;
      RECT 79.555000  23.335000 80.115000  23.405000 ;
      RECT 79.605000  17.275000 80.000000  19.205000 ;
      RECT 79.605000  21.045000 80.115000  21.115000 ;
      RECT 79.605000  31.795000 80.115000  31.865000 ;
      RECT 79.605000  33.975000 80.115000  34.045000 ;
      RECT 79.625000  23.405000 80.115000  23.475000 ;
      RECT 79.675000  20.975000 80.115000  21.045000 ;
      RECT 79.675000  31.725000 80.115000  31.795000 ;
      RECT 79.675000  34.045000 80.115000  34.115000 ;
      RECT 79.695000  23.475000 80.115000  23.545000 ;
      RECT 79.745000  20.905000 80.115000  20.975000 ;
      RECT 79.745000  31.655000 80.115000  31.725000 ;
      RECT 79.745000  34.115000 80.115000  34.185000 ;
      RECT 79.765000  23.545000 80.115000  23.615000 ;
      RECT 79.815000  20.835000 80.115000  20.905000 ;
      RECT 79.815000  31.585000 80.115000  31.655000 ;
      RECT 79.815000  34.185000 80.115000  34.255000 ;
      RECT 79.835000  23.615000 80.115000  23.685000 ;
      RECT 79.885000  19.485000 80.115000  20.765000 ;
      RECT 79.885000  20.765000 80.115000  20.835000 ;
      RECT 79.885000  23.685000 80.115000  23.735000 ;
      RECT 79.885000  23.735000 80.115000  25.015000 ;
      RECT 79.885000  30.120000 80.115000  31.515000 ;
      RECT 79.885000  31.515000 80.115000  31.585000 ;
      RECT 79.885000  34.255000 80.115000  34.325000 ;
      RECT 79.885000  34.325000 80.115000  35.725000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  3.095000   4.591000 ;
      RECT  0.000000   0.000000  3.235000   4.533000 ;
      RECT  0.000000   4.533000  3.942000   5.240000 ;
      RECT  0.000000   4.591000  3.095000   4.660000 ;
      RECT  0.000000   4.591000  3.095000   4.660000 ;
      RECT  0.000000   4.660000  3.164000   4.730000 ;
      RECT  0.000000   4.660000  3.164000   4.730000 ;
      RECT  0.000000   4.730000  3.234000   4.800000 ;
      RECT  0.000000   4.730000  3.234000   4.800000 ;
      RECT  0.000000   4.800000  3.304000   4.870000 ;
      RECT  0.000000   4.800000  3.304000   4.870000 ;
      RECT  0.000000   4.870000  3.374000   4.940000 ;
      RECT  0.000000   4.870000  3.374000   4.940000 ;
      RECT  0.000000   4.940000  3.444000   5.010000 ;
      RECT  0.000000   4.940000  3.444000   5.010000 ;
      RECT  0.000000   5.010000  3.514000   5.080000 ;
      RECT  0.000000   5.010000  3.514000   5.080000 ;
      RECT  0.000000   5.080000  3.584000   5.150000 ;
      RECT  0.000000   5.080000  3.584000   5.150000 ;
      RECT  0.000000   5.150000  3.654000   5.220000 ;
      RECT  0.000000   5.150000  3.654000   5.220000 ;
      RECT  0.000000   5.220000  3.724000   5.290000 ;
      RECT  0.000000   5.220000  3.724000   5.290000 ;
      RECT  0.000000   5.240000  5.260000   5.433000 ;
      RECT  0.000000   5.290000  3.794000   5.360000 ;
      RECT  0.000000   5.290000  3.794000   5.360000 ;
      RECT  0.000000   5.360000  3.864000   5.380000 ;
      RECT  0.000000   5.360000  3.864000   5.380000 ;
      RECT  0.000000   5.380000  5.009000   5.435000 ;
      RECT  0.000000   5.380000  5.009000   5.435000 ;
      RECT  0.000000   5.433000  5.260000   8.408000 ;
      RECT  0.000000   5.435000  5.064000   5.490000 ;
      RECT  0.000000   5.435000  5.064000   5.490000 ;
      RECT  0.000000   5.491000  5.120000   8.496000 ;
      RECT  0.000000   8.408000  6.435000   9.583000 ;
      RECT  0.000000   8.466000  5.120000   8.535000 ;
      RECT  0.000000   8.466000  5.120000   8.535000 ;
      RECT  0.000000   8.535000  5.189000   8.605000 ;
      RECT  0.000000   8.535000  5.189000   8.605000 ;
      RECT  0.000000   8.605000  5.259000   8.675000 ;
      RECT  0.000000   8.605000  5.259000   8.675000 ;
      RECT  0.000000   8.675000  5.329000   8.745000 ;
      RECT  0.000000   8.675000  5.329000   8.745000 ;
      RECT  0.000000   8.745000  5.399000   8.815000 ;
      RECT  0.000000   8.745000  5.399000   8.815000 ;
      RECT  0.000000   8.815000  5.469000   8.885000 ;
      RECT  0.000000   8.815000  5.469000   8.885000 ;
      RECT  0.000000   8.885000  5.539000   8.955000 ;
      RECT  0.000000   8.885000  5.539000   8.955000 ;
      RECT  0.000000   8.955000  5.609000   9.025000 ;
      RECT  0.000000   8.955000  5.609000   9.025000 ;
      RECT  0.000000   9.025000  5.679000   9.095000 ;
      RECT  0.000000   9.025000  5.679000   9.095000 ;
      RECT  0.000000   9.095000  5.749000   9.165000 ;
      RECT  0.000000   9.095000  5.749000   9.165000 ;
      RECT  0.000000   9.165000  5.819000   9.235000 ;
      RECT  0.000000   9.165000  5.819000   9.235000 ;
      RECT  0.000000   9.235000  5.889000   9.305000 ;
      RECT  0.000000   9.235000  5.889000   9.305000 ;
      RECT  0.000000   9.305000  5.959000   9.375000 ;
      RECT  0.000000   9.305000  5.959000   9.375000 ;
      RECT  0.000000   9.375000  6.029000   9.445000 ;
      RECT  0.000000   9.375000  6.029000   9.445000 ;
      RECT  0.000000   9.445000  6.099000   9.515000 ;
      RECT  0.000000   9.445000  6.099000   9.515000 ;
      RECT  0.000000   9.515000  6.169000   9.585000 ;
      RECT  0.000000   9.515000  6.169000   9.585000 ;
      RECT  0.000000   9.583000  6.435000  38.762000 ;
      RECT  0.000000   9.585000  6.239000   9.640000 ;
      RECT  0.000000   9.585000  6.239000   9.640000 ;
      RECT  0.000000   9.641000  6.295000  38.704000 ;
      RECT  0.000000  38.704000  6.224000  38.775000 ;
      RECT  0.000000  38.704000  6.224000  38.775000 ;
      RECT  0.000000  38.762000  5.835000  39.362000 ;
      RECT  0.000000  38.775000  6.154000  38.845000 ;
      RECT  0.000000  38.775000  6.154000  38.845000 ;
      RECT  0.000000  38.845000  6.084000  38.915000 ;
      RECT  0.000000  38.845000  6.084000  38.915000 ;
      RECT  0.000000  38.915000  6.014000  38.985000 ;
      RECT  0.000000  38.915000  6.014000  38.985000 ;
      RECT  0.000000  38.985000  5.944000  39.055000 ;
      RECT  0.000000  38.985000  5.944000  39.055000 ;
      RECT  0.000000  39.055000  5.874000  39.125000 ;
      RECT  0.000000  39.055000  5.874000  39.125000 ;
      RECT  0.000000  39.125000  5.804000  39.195000 ;
      RECT  0.000000  39.125000  5.804000  39.195000 ;
      RECT  0.000000  39.195000  5.734000  39.265000 ;
      RECT  0.000000  39.195000  5.734000  39.265000 ;
      RECT  0.000000  39.265000  5.694000  39.305000 ;
      RECT  0.000000  39.265000  5.694000  39.305000 ;
      RECT  0.000000  39.304000  5.685000  53.624000 ;
      RECT  0.000000  39.304000  5.695000  42.859000 ;
      RECT  0.000000  39.362000  5.835000  42.917000 ;
      RECT  0.000000  42.859000  5.689000  42.865000 ;
      RECT  0.000000  42.859000  5.689000  42.865000 ;
      RECT  0.000000  42.865000  5.684000  42.870000 ;
      RECT  0.000000  42.865000  5.684000  42.870000 ;
      RECT  0.000000  42.869000  5.685000  43.905000 ;
      RECT  0.000000  42.917000  5.825000  42.927000 ;
      RECT  0.000000  42.927000  5.825000  43.765000 ;
      RECT  0.000000  43.765000  8.055000  44.017000 ;
      RECT  0.000000  43.905000  7.915000  53.624000 ;
      RECT  0.000000  43.905000  7.944000  43.930000 ;
      RECT  0.000000  43.905000  7.944000  43.930000 ;
      RECT  0.000000  43.930000  7.919000  43.955000 ;
      RECT  0.000000  43.930000  7.919000  43.955000 ;
      RECT  0.000000  43.955000  7.914000  43.960000 ;
      RECT  0.000000  43.955000  7.914000  43.960000 ;
      RECT  0.000000  43.959000  7.915000  53.624000 ;
      RECT  0.000000  44.017000  8.055000  53.682000 ;
      RECT  0.000000  53.624000  7.844000  53.695000 ;
      RECT  0.000000  53.624000  7.844000  53.695000 ;
      RECT  0.000000  53.682000  7.835000  53.902000 ;
      RECT  0.000000  53.695000  7.774000  53.765000 ;
      RECT  0.000000  53.695000  7.774000  53.765000 ;
      RECT  0.000000  53.765000  7.704000  53.835000 ;
      RECT  0.000000  53.765000  7.704000  53.835000 ;
      RECT  0.000000  53.835000  7.694000  53.845000 ;
      RECT  0.000000  53.835000  7.694000  53.845000 ;
      RECT  0.000000  53.844000  7.695000  55.684000 ;
      RECT  0.000000  53.902000  7.835000  55.742000 ;
      RECT  0.000000  55.684000  7.035000  73.841000 ;
      RECT  0.000000  55.684000  7.035000  73.841000 ;
      RECT  0.000000  55.684000  7.035000  73.841000 ;
      RECT  0.000000  55.684000  7.035000  73.841000 ;
      RECT  0.000000  55.684000  7.624000  55.755000 ;
      RECT  0.000000  55.684000  7.624000  55.755000 ;
      RECT  0.000000  55.742000  7.175000  56.402000 ;
      RECT  0.000000  55.755000  7.554000  55.825000 ;
      RECT  0.000000  55.755000  7.554000  55.825000 ;
      RECT  0.000000  55.825000  7.484000  55.895000 ;
      RECT  0.000000  55.825000  7.484000  55.895000 ;
      RECT  0.000000  55.895000  7.414000  55.965000 ;
      RECT  0.000000  55.895000  7.414000  55.965000 ;
      RECT  0.000000  55.965000  7.344000  56.035000 ;
      RECT  0.000000  55.965000  7.344000  56.035000 ;
      RECT  0.000000  56.035000  7.274000  56.105000 ;
      RECT  0.000000  56.035000  7.274000  56.105000 ;
      RECT  0.000000  56.105000  7.204000  56.175000 ;
      RECT  0.000000  56.105000  7.204000  56.175000 ;
      RECT  0.000000  56.175000  7.134000  56.245000 ;
      RECT  0.000000  56.175000  7.134000  56.245000 ;
      RECT  0.000000  56.245000  7.064000  56.315000 ;
      RECT  0.000000  56.245000  7.064000  56.315000 ;
      RECT  0.000000  56.315000  7.034000  56.345000 ;
      RECT  0.000000  56.315000  7.034000  56.345000 ;
      RECT  0.000000  56.402000  7.175000  73.783000 ;
      RECT  0.000000  73.783000  7.665000  74.273000 ;
      RECT  0.000000  73.841000  7.035000  73.910000 ;
      RECT  0.000000  73.841000  7.035000  73.910000 ;
      RECT  0.000000  73.910000  7.104000  73.980000 ;
      RECT  0.000000  73.910000  7.104000  73.980000 ;
      RECT  0.000000  73.980000  7.174000  74.050000 ;
      RECT  0.000000  73.980000  7.174000  74.050000 ;
      RECT  0.000000  74.050000  7.244000  74.120000 ;
      RECT  0.000000  74.050000  7.244000  74.120000 ;
      RECT  0.000000  74.120000  7.314000  74.190000 ;
      RECT  0.000000  74.120000  7.314000  74.190000 ;
      RECT  0.000000  74.190000  7.384000  74.260000 ;
      RECT  0.000000  74.190000  7.384000  74.260000 ;
      RECT  0.000000  74.260000  7.454000  74.330000 ;
      RECT  0.000000  74.260000  7.454000  74.330000 ;
      RECT  0.000000  74.273000  7.665000  74.848000 ;
      RECT  0.000000  74.331000  7.525000  74.906000 ;
      RECT  0.000000  74.848000  8.070000  75.253000 ;
      RECT  0.000000  74.906000  7.525000  74.965000 ;
      RECT  0.000000  74.906000  7.525000  74.965000 ;
      RECT  0.000000  74.906000  7.525000  74.975000 ;
      RECT  0.000000  74.965000  7.584000  75.020000 ;
      RECT  0.000000  74.965000  7.584000  75.020000 ;
      RECT  0.000000  74.975000  7.594000  75.045000 ;
      RECT  0.000000  75.021000  7.640000  75.311000 ;
      RECT  0.000000  75.045000  7.664000  75.115000 ;
      RECT  0.000000  75.115000  7.734000  75.185000 ;
      RECT  0.000000  75.185000  7.804000  75.255000 ;
      RECT  0.000000  75.253000  8.070000  77.057000 ;
      RECT  0.000000  75.255000  7.874000  75.310000 ;
      RECT  0.000000  75.311000  7.930000  77.005000 ;
      RECT  0.000000  77.005000  7.640000  78.316000 ;
      RECT  0.000000  77.057000  7.982000  77.145000 ;
      RECT  0.000000  77.145000  7.780000  77.685000 ;
      RECT  0.000000  77.685000 76.775000  96.137000 ;
      RECT  0.000000  77.825000 76.635000  96.079000 ;
      RECT  0.000000  96.079000 76.564000  96.150000 ;
      RECT  0.000000  96.079000 76.564000  96.150000 ;
      RECT  0.000000  96.137000 76.547000  96.365000 ;
      RECT  0.000000  96.150000 76.494000  96.220000 ;
      RECT  0.000000  96.150000 76.494000  96.220000 ;
      RECT  0.000000  96.220000 76.424000  96.290000 ;
      RECT  0.000000  96.220000 76.424000  96.290000 ;
      RECT  0.000000  96.290000 76.354000  96.360000 ;
      RECT  0.000000  96.290000 76.354000  96.360000 ;
      RECT  0.000000  96.360000 76.284000  96.430000 ;
      RECT  0.000000  96.360000 76.284000  96.430000 ;
      RECT  0.000000  96.365000 80.000000 106.585000 ;
      RECT  0.000000  96.430000 76.214000  96.500000 ;
      RECT  0.000000  96.430000 76.214000  96.500000 ;
      RECT  0.000000  96.500000 76.209000  96.505000 ;
      RECT  0.000000  96.500000 76.209000  96.505000 ;
      RECT  0.000000  96.505000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.740000 106.585000 80.000000 118.955000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  3.745000   0.000000  5.280000   4.317000 ;
      RECT  3.745000   4.317000  5.280000   4.533000 ;
      RECT  3.885000   0.000000  5.140000   4.259000 ;
      RECT  3.956000   4.259000  5.140000   4.330000 ;
      RECT  3.961000   4.533000  5.477000   4.730000 ;
      RECT  4.026000   4.330000  5.140000   4.400000 ;
      RECT  4.096000   4.400000  5.140000   4.470000 ;
      RECT  4.166000   4.470000  5.140000   4.540000 ;
      RECT  4.216000   4.540000  5.140000   4.590000 ;
      RECT  5.283000   4.730000  5.964000   5.217000 ;
      RECT  5.770000   5.217000  6.180000   5.433000 ;
      RECT  5.770000   5.433000  6.180000   6.192000 ;
      RECT  5.770000   6.192000  6.087000   6.285000 ;
      RECT  5.770000   6.825000  8.305000   6.920000 ;
      RECT  5.770000   6.920000 13.830000   8.192000 ;
      RECT  5.770000   8.192000 13.830000   9.367000 ;
      RECT  5.790000   0.000000  5.990000   1.608000 ;
      RECT  5.790000   1.608000  8.305000   3.923000 ;
      RECT  5.790000   3.923000  8.305000   4.317000 ;
      RECT  5.790000   4.317000  8.305000   5.217000 ;
      RECT  5.845000   2.335000  6.519000   2.405000 ;
      RECT  5.845000   2.405000  6.589000   2.475000 ;
      RECT  5.845000   2.475000  6.659000   2.545000 ;
      RECT  5.845000   2.545000  6.729000   2.595000 ;
      RECT  5.885000   2.595000  6.779000   2.635000 ;
      RECT  5.910000   6.965000  8.165000   7.060000 ;
      RECT  5.910000   7.060000 13.690000   7.344000 ;
      RECT  5.910000   7.344000 13.690000   8.134000 ;
      RECT  5.925000   2.635000  6.819000   2.675000 ;
      RECT  5.930000   1.815000  5.999000   1.885000 ;
      RECT  5.930000   1.885000  6.069000   1.955000 ;
      RECT  5.930000   1.955000  6.139000   2.025000 ;
      RECT  5.930000   2.025000  6.209000   2.095000 ;
      RECT  5.930000   2.095000  6.279000   2.165000 ;
      RECT  5.930000   2.165000  6.349000   2.235000 ;
      RECT  5.930000   2.235000  6.419000   2.305000 ;
      RECT  5.930000   2.305000  6.489000   2.335000 ;
      RECT  5.930000   2.675000  6.859000   2.680000 ;
      RECT  5.930000   2.680000  6.864000   2.750000 ;
      RECT  5.930000   2.750000  6.934000   2.820000 ;
      RECT  5.930000   2.820000  7.004000   2.890000 ;
      RECT  5.930000   2.890000  7.074000   2.960000 ;
      RECT  5.930000   2.960000  7.144000   3.030000 ;
      RECT  5.930000   3.030000  7.214000   3.100000 ;
      RECT  5.930000   3.100000  7.284000   3.170000 ;
      RECT  5.930000   3.170000  7.354000   3.240000 ;
      RECT  5.930000   3.240000  7.424000   3.310000 ;
      RECT  5.930000   3.310000  7.494000   3.380000 ;
      RECT  5.930000   3.380000  7.564000   3.450000 ;
      RECT  5.930000   3.450000  7.634000   3.520000 ;
      RECT  5.930000   3.520000  7.704000   3.590000 ;
      RECT  5.930000   3.590000  7.774000   3.660000 ;
      RECT  5.930000   3.660000  7.844000   3.730000 ;
      RECT  5.930000   3.730000  7.914000   3.800000 ;
      RECT  5.930000   3.800000  7.984000   3.870000 ;
      RECT  5.930000   3.870000  8.054000   3.940000 ;
      RECT  5.930000   3.940000  8.124000   3.980000 ;
      RECT  5.930000   3.981000  8.165000   4.259000 ;
      RECT  5.981000   8.134000 13.690000   8.205000 ;
      RECT  5.981000   8.134000 13.690000   8.205000 ;
      RECT  6.001000   4.259000  8.165000   4.330000 ;
      RECT  6.051000   8.205000 13.690000   8.275000 ;
      RECT  6.051000   8.205000 13.690000   8.275000 ;
      RECT  6.071000   4.330000  8.165000   4.400000 ;
      RECT  6.121000   8.275000 13.690000   8.345000 ;
      RECT  6.121000   8.275000 13.690000   8.345000 ;
      RECT  6.141000   4.400000  8.165000   4.470000 ;
      RECT  6.191000   8.345000 13.690000   8.415000 ;
      RECT  6.191000   8.345000 13.690000   8.415000 ;
      RECT  6.211000   4.470000  8.165000   4.540000 ;
      RECT  6.261000   8.415000 13.690000   8.485000 ;
      RECT  6.261000   8.415000 13.690000   8.485000 ;
      RECT  6.281000   4.540000  8.165000   4.610000 ;
      RECT  6.331000   8.485000 13.690000   8.555000 ;
      RECT  6.331000   8.485000 13.690000   8.555000 ;
      RECT  6.345000  39.578000  9.165000  42.907000 ;
      RECT  6.345000  42.907000  9.145000  42.927000 ;
      RECT  6.351000   4.610000  8.165000   4.680000 ;
      RECT  6.365000  42.927000  8.307000  43.765000 ;
      RECT  6.401000   8.555000 13.690000   8.625000 ;
      RECT  6.401000   8.555000 13.690000   8.625000 ;
      RECT  6.421000   4.680000  8.165000   4.750000 ;
      RECT  6.471000   8.625000 13.690000   8.695000 ;
      RECT  6.471000   8.625000 13.690000   8.695000 ;
      RECT  6.485000  39.636000 12.169000  39.705000 ;
      RECT  6.485000  39.636000 12.169000  39.705000 ;
      RECT  6.485000  39.705000 12.099000  39.775000 ;
      RECT  6.485000  39.705000 12.099000  39.775000 ;
      RECT  6.485000  39.775000 12.029000  39.845000 ;
      RECT  6.485000  39.775000 12.029000  39.845000 ;
      RECT  6.485000  39.845000 11.959000  39.915000 ;
      RECT  6.485000  39.845000 11.959000  39.915000 ;
      RECT  6.485000  39.915000 11.889000  39.985000 ;
      RECT  6.485000  39.915000 11.889000  39.985000 ;
      RECT  6.485000  39.985000 11.819000  40.055000 ;
      RECT  6.485000  39.985000 11.819000  40.055000 ;
      RECT  6.485000  40.055000 11.749000  40.125000 ;
      RECT  6.485000  40.055000 11.749000  40.125000 ;
      RECT  6.485000  40.125000 11.679000  40.195000 ;
      RECT  6.485000  40.125000 11.679000  40.195000 ;
      RECT  6.485000  40.195000 11.609000  40.265000 ;
      RECT  6.485000  40.195000 11.609000  40.265000 ;
      RECT  6.485000  40.265000 11.539000  40.335000 ;
      RECT  6.485000  40.265000 11.539000  40.335000 ;
      RECT  6.485000  40.335000 11.469000  40.405000 ;
      RECT  6.485000  40.335000 11.469000  40.405000 ;
      RECT  6.485000  40.405000 11.399000  40.475000 ;
      RECT  6.485000  40.405000 11.399000  40.475000 ;
      RECT  6.485000  40.475000 11.329000  40.545000 ;
      RECT  6.485000  40.475000 11.329000  40.545000 ;
      RECT  6.485000  40.545000 11.259000  40.615000 ;
      RECT  6.485000  40.545000 11.259000  40.615000 ;
      RECT  6.485000  40.615000 11.189000  40.685000 ;
      RECT  6.485000  40.615000 11.189000  40.685000 ;
      RECT  6.485000  40.685000 11.119000  40.755000 ;
      RECT  6.485000  40.685000 11.119000  40.755000 ;
      RECT  6.485000  40.755000 11.049000  40.825000 ;
      RECT  6.485000  40.755000 11.049000  40.825000 ;
      RECT  6.485000  40.825000 10.979000  40.895000 ;
      RECT  6.485000  40.825000 10.979000  40.895000 ;
      RECT  6.485000  40.895000 10.909000  40.965000 ;
      RECT  6.485000  40.895000 10.909000  40.965000 ;
      RECT  6.485000  40.965000 10.839000  41.035000 ;
      RECT  6.485000  40.965000 10.839000  41.035000 ;
      RECT  6.485000  41.035000 10.769000  41.105000 ;
      RECT  6.485000  41.035000 10.769000  41.105000 ;
      RECT  6.485000  41.105000 10.699000  41.175000 ;
      RECT  6.485000  41.105000 10.699000  41.175000 ;
      RECT  6.485000  41.175000 10.629000  41.245000 ;
      RECT  6.485000  41.175000 10.629000  41.245000 ;
      RECT  6.485000  41.245000 10.559000  41.315000 ;
      RECT  6.485000  41.245000 10.559000  41.315000 ;
      RECT  6.485000  41.315000 10.489000  41.385000 ;
      RECT  6.485000  41.315000 10.489000  41.385000 ;
      RECT  6.485000  41.385000 10.419000  41.455000 ;
      RECT  6.485000  41.385000 10.419000  41.455000 ;
      RECT  6.485000  41.455000 10.349000  41.525000 ;
      RECT  6.485000  41.455000 10.349000  41.525000 ;
      RECT  6.485000  41.525000 10.279000  41.595000 ;
      RECT  6.485000  41.525000 10.279000  41.595000 ;
      RECT  6.485000  41.595000 10.209000  41.665000 ;
      RECT  6.485000  41.595000 10.209000  41.665000 ;
      RECT  6.485000  41.665000 10.139000  41.735000 ;
      RECT  6.485000  41.665000 10.139000  41.735000 ;
      RECT  6.485000  41.735000 10.069000  41.805000 ;
      RECT  6.485000  41.735000 10.069000  41.805000 ;
      RECT  6.485000  41.805000  9.999000  41.875000 ;
      RECT  6.485000  41.805000  9.999000  41.875000 ;
      RECT  6.485000  41.875000  9.929000  41.945000 ;
      RECT  6.485000  41.875000  9.929000  41.945000 ;
      RECT  6.485000  41.945000  9.859000  42.015000 ;
      RECT  6.485000  41.945000  9.859000  42.015000 ;
      RECT  6.485000  42.015000  9.789000  42.085000 ;
      RECT  6.485000  42.015000  9.789000  42.085000 ;
      RECT  6.485000  42.085000  9.719000  42.155000 ;
      RECT  6.485000  42.085000  9.719000  42.155000 ;
      RECT  6.485000  42.155000  9.649000  42.225000 ;
      RECT  6.485000  42.155000  9.649000  42.225000 ;
      RECT  6.485000  42.225000  9.579000  42.295000 ;
      RECT  6.485000  42.225000  9.579000  42.295000 ;
      RECT  6.485000  42.295000  9.509000  42.365000 ;
      RECT  6.485000  42.295000  9.509000  42.365000 ;
      RECT  6.485000  42.365000  9.439000  42.435000 ;
      RECT  6.485000  42.365000  9.439000  42.435000 ;
      RECT  6.485000  42.435000  9.369000  42.505000 ;
      RECT  6.485000  42.435000  9.369000  42.505000 ;
      RECT  6.485000  42.505000  9.299000  42.575000 ;
      RECT  6.485000  42.505000  9.299000  42.575000 ;
      RECT  6.485000  42.575000  9.229000  42.645000 ;
      RECT  6.485000  42.575000  9.229000  42.645000 ;
      RECT  6.485000  42.645000  9.159000  42.715000 ;
      RECT  6.485000  42.645000  9.159000  42.715000 ;
      RECT  6.485000  42.715000  9.089000  42.785000 ;
      RECT  6.485000  42.715000  9.089000  42.785000 ;
      RECT  6.485000  42.785000  9.024000  42.850000 ;
      RECT  6.485000  42.785000  9.024000  42.850000 ;
      RECT  6.491000   4.750000  8.165000   4.820000 ;
      RECT  6.496000  42.849000  9.014000  42.860000 ;
      RECT  6.496000  42.849000  9.014000  42.860000 ;
      RECT  6.505000  42.869000  8.934000  42.940000 ;
      RECT  6.505000  42.869000  8.934000  42.940000 ;
      RECT  6.505000  42.940000  8.864000  43.010000 ;
      RECT  6.505000  42.940000  8.864000  43.010000 ;
      RECT  6.505000  43.010000  8.794000  43.080000 ;
      RECT  6.505000  43.010000  8.794000  43.080000 ;
      RECT  6.505000  43.080000  8.724000  43.150000 ;
      RECT  6.505000  43.080000  8.724000  43.150000 ;
      RECT  6.505000  43.150000  8.654000  43.220000 ;
      RECT  6.505000  43.150000  8.654000  43.220000 ;
      RECT  6.505000  43.220000  8.584000  43.290000 ;
      RECT  6.505000  43.220000  8.584000  43.290000 ;
      RECT  6.505000  43.290000  8.514000  43.360000 ;
      RECT  6.505000  43.290000  8.514000  43.360000 ;
      RECT  6.505000  43.360000  8.444000  43.430000 ;
      RECT  6.505000  43.360000  8.444000  43.430000 ;
      RECT  6.505000  43.430000  8.374000  43.500000 ;
      RECT  6.505000  43.430000  8.374000  43.500000 ;
      RECT  6.505000  43.500000  8.304000  43.570000 ;
      RECT  6.505000  43.500000  8.304000  43.570000 ;
      RECT  6.505000  43.570000  8.234000  43.640000 ;
      RECT  6.505000  43.570000  8.234000  43.640000 ;
      RECT  6.505000  43.640000  8.164000  43.710000 ;
      RECT  6.505000  43.640000  8.164000  43.710000 ;
      RECT  6.505000  43.710000  8.094000  43.780000 ;
      RECT  6.505000  43.710000  8.094000  43.780000 ;
      RECT  6.505000  43.780000  8.024000  43.850000 ;
      RECT  6.505000  43.780000  8.024000  43.850000 ;
      RECT  6.505000  43.850000  7.969000  43.905000 ;
      RECT  6.505000  43.850000  7.969000  43.905000 ;
      RECT  6.506000  42.860000  9.004000  42.870000 ;
      RECT  6.506000  42.860000  9.004000  42.870000 ;
      RECT  6.526000  39.595000 12.239000  39.635000 ;
      RECT  6.526000  39.595000 12.239000  39.635000 ;
      RECT  6.530000   0.000000 12.615000   1.382000 ;
      RECT  6.530000   1.382000 12.615000   3.697000 ;
      RECT  6.541000   8.695000 13.690000   8.765000 ;
      RECT  6.541000   8.695000 13.690000   8.765000 ;
      RECT  6.561000   4.820000  8.165000   4.890000 ;
      RECT  6.596000  39.525000 12.279000  39.595000 ;
      RECT  6.596000  39.525000 12.279000  39.595000 ;
      RECT  6.611000   8.765000 13.690000   8.835000 ;
      RECT  6.611000   8.765000 13.690000   8.835000 ;
      RECT  6.631000   4.890000  8.165000   4.960000 ;
      RECT  6.666000  39.455000 12.349000  39.525000 ;
      RECT  6.666000  39.455000 12.349000  39.525000 ;
      RECT  6.670000   0.000000 12.475000   1.324000 ;
      RECT  6.681000   8.835000 13.690000   8.905000 ;
      RECT  6.681000   8.835000 13.690000   8.905000 ;
      RECT  6.690000   5.217000  8.305000   6.825000 ;
      RECT  6.701000   4.960000  8.165000   5.030000 ;
      RECT  6.736000  39.385000 12.419000  39.455000 ;
      RECT  6.736000  39.385000 12.419000  39.455000 ;
      RECT  6.741000   1.324000 12.475000   1.395000 ;
      RECT  6.741000   1.324000 12.475000   1.395000 ;
      RECT  6.751000   8.905000 13.690000   8.975000 ;
      RECT  6.751000   8.905000 13.690000   8.975000 ;
      RECT  6.771000   5.030000  8.165000   5.100000 ;
      RECT  6.806000  39.315000 12.489000  39.385000 ;
      RECT  6.806000  39.315000 12.489000  39.385000 ;
      RECT  6.811000   1.395000 12.475000   1.465000 ;
      RECT  6.811000   1.395000 12.475000   1.465000 ;
      RECT  6.821000   8.975000 13.690000   9.045000 ;
      RECT  6.821000   8.975000 13.690000   9.045000 ;
      RECT  6.830000   5.159000  8.165000   6.965000 ;
      RECT  6.831000   5.100000  8.165000   5.160000 ;
      RECT  6.876000  39.245000 12.559000  39.315000 ;
      RECT  6.876000  39.245000 12.559000  39.315000 ;
      RECT  6.881000   1.465000 12.475000   1.535000 ;
      RECT  6.881000   1.465000 12.475000   1.535000 ;
      RECT  6.891000   9.045000 13.690000   9.115000 ;
      RECT  6.891000   9.045000 13.690000   9.115000 ;
      RECT  6.945000   9.367000 13.830000  18.283000 ;
      RECT  6.945000  18.283000 15.245000  19.698000 ;
      RECT  6.945000  19.698000 15.245000  31.487000 ;
      RECT  6.945000  31.487000 14.830000  31.902000 ;
      RECT  6.945000  31.902000 14.830000  37.242000 ;
      RECT  6.945000  37.242000 13.094000  38.978000 ;
      RECT  6.945000  38.978000 12.494000  39.578000 ;
      RECT  6.946000  39.175000 12.629000  39.245000 ;
      RECT  6.946000  39.175000 12.629000  39.245000 ;
      RECT  6.951000   1.535000 12.475000   1.605000 ;
      RECT  6.951000   1.535000 12.475000   1.605000 ;
      RECT  6.961000   9.115000 13.690000   9.185000 ;
      RECT  6.961000   9.115000 13.690000   9.185000 ;
      RECT  7.016000  39.105000 12.699000  39.175000 ;
      RECT  7.016000  39.105000 12.699000  39.175000 ;
      RECT  7.021000   1.605000 12.475000   1.675000 ;
      RECT  7.021000   1.605000 12.475000   1.675000 ;
      RECT  7.031000   9.185000 13.690000   9.255000 ;
      RECT  7.031000   9.185000 13.690000   9.255000 ;
      RECT  7.085000   9.309000 13.690000  18.341000 ;
      RECT  7.085000  18.341000 13.690000  18.410000 ;
      RECT  7.085000  18.341000 13.690000  18.410000 ;
      RECT  7.085000  18.410000 13.759000  18.480000 ;
      RECT  7.085000  18.410000 13.759000  18.480000 ;
      RECT  7.085000  18.480000 13.829000  18.550000 ;
      RECT  7.085000  18.480000 13.829000  18.550000 ;
      RECT  7.085000  18.550000 13.899000  18.620000 ;
      RECT  7.085000  18.550000 13.899000  18.620000 ;
      RECT  7.085000  18.620000 13.969000  18.690000 ;
      RECT  7.085000  18.620000 13.969000  18.690000 ;
      RECT  7.085000  18.690000 14.039000  18.760000 ;
      RECT  7.085000  18.690000 14.039000  18.760000 ;
      RECT  7.085000  18.760000 14.109000  18.830000 ;
      RECT  7.085000  18.760000 14.109000  18.830000 ;
      RECT  7.085000  18.830000 14.179000  18.900000 ;
      RECT  7.085000  18.830000 14.179000  18.900000 ;
      RECT  7.085000  18.900000 14.249000  18.970000 ;
      RECT  7.085000  18.900000 14.249000  18.970000 ;
      RECT  7.085000  18.970000 14.319000  19.040000 ;
      RECT  7.085000  18.970000 14.319000  19.040000 ;
      RECT  7.085000  19.040000 14.389000  19.110000 ;
      RECT  7.085000  19.040000 14.389000  19.110000 ;
      RECT  7.085000  19.110000 14.459000  19.180000 ;
      RECT  7.085000  19.110000 14.459000  19.180000 ;
      RECT  7.085000  19.180000 14.529000  19.250000 ;
      RECT  7.085000  19.180000 14.529000  19.250000 ;
      RECT  7.085000  19.250000 14.599000  19.320000 ;
      RECT  7.085000  19.250000 14.599000  19.320000 ;
      RECT  7.085000  19.320000 14.669000  19.390000 ;
      RECT  7.085000  19.320000 14.669000  19.390000 ;
      RECT  7.085000  19.390000 14.739000  19.460000 ;
      RECT  7.085000  19.390000 14.739000  19.460000 ;
      RECT  7.085000  19.460000 14.809000  19.530000 ;
      RECT  7.085000  19.460000 14.809000  19.530000 ;
      RECT  7.085000  19.530000 14.879000  19.600000 ;
      RECT  7.085000  19.530000 14.879000  19.600000 ;
      RECT  7.085000  19.600000 14.949000  19.670000 ;
      RECT  7.085000  19.600000 14.949000  19.670000 ;
      RECT  7.085000  19.670000 15.019000  19.740000 ;
      RECT  7.085000  19.670000 15.019000  19.740000 ;
      RECT  7.085000  19.740000 15.089000  19.755000 ;
      RECT  7.085000  19.740000 15.089000  19.755000 ;
      RECT  7.085000  19.756000 15.105000  31.429000 ;
      RECT  7.085000  31.429000 15.034000  31.500000 ;
      RECT  7.085000  31.429000 15.034000  31.500000 ;
      RECT  7.085000  31.500000 14.964000  31.570000 ;
      RECT  7.085000  31.500000 14.964000  31.570000 ;
      RECT  7.085000  31.570000 14.894000  31.640000 ;
      RECT  7.085000  31.570000 14.894000  31.640000 ;
      RECT  7.085000  31.640000 14.824000  31.710000 ;
      RECT  7.085000  31.640000 14.824000  31.710000 ;
      RECT  7.085000  31.710000 14.754000  31.780000 ;
      RECT  7.085000  31.710000 14.754000  31.780000 ;
      RECT  7.085000  31.780000 14.689000  31.845000 ;
      RECT  7.085000  31.780000 14.689000  31.845000 ;
      RECT  7.085000  31.844000 14.690000  37.184000 ;
      RECT  7.085000  37.184000 14.619000  37.255000 ;
      RECT  7.085000  37.184000 14.619000  37.255000 ;
      RECT  7.085000  37.255000 14.549000  37.325000 ;
      RECT  7.085000  37.255000 14.549000  37.325000 ;
      RECT  7.085000  37.325000 14.479000  37.395000 ;
      RECT  7.085000  37.325000 14.479000  37.395000 ;
      RECT  7.085000  37.395000 14.409000  37.465000 ;
      RECT  7.085000  37.395000 14.409000  37.465000 ;
      RECT  7.085000  37.465000 14.339000  37.535000 ;
      RECT  7.085000  37.465000 14.339000  37.535000 ;
      RECT  7.085000  37.535000 14.269000  37.605000 ;
      RECT  7.085000  37.535000 14.269000  37.605000 ;
      RECT  7.085000  37.605000 14.199000  37.675000 ;
      RECT  7.085000  37.605000 14.199000  37.675000 ;
      RECT  7.085000  37.675000 14.129000  37.745000 ;
      RECT  7.085000  37.675000 14.129000  37.745000 ;
      RECT  7.085000  37.745000 14.059000  37.815000 ;
      RECT  7.085000  37.745000 14.059000  37.815000 ;
      RECT  7.085000  37.815000 13.989000  37.885000 ;
      RECT  7.085000  37.815000 13.989000  37.885000 ;
      RECT  7.085000  37.885000 13.919000  37.955000 ;
      RECT  7.085000  37.885000 13.919000  37.955000 ;
      RECT  7.085000  37.955000 13.849000  38.025000 ;
      RECT  7.085000  37.955000 13.849000  38.025000 ;
      RECT  7.085000  38.025000 13.779000  38.095000 ;
      RECT  7.085000  38.025000 13.779000  38.095000 ;
      RECT  7.085000  38.095000 13.709000  38.165000 ;
      RECT  7.085000  38.095000 13.709000  38.165000 ;
      RECT  7.085000  38.165000 13.639000  38.235000 ;
      RECT  7.085000  38.165000 13.639000  38.235000 ;
      RECT  7.085000  38.235000 13.569000  38.305000 ;
      RECT  7.085000  38.235000 13.569000  38.305000 ;
      RECT  7.085000  38.305000 13.499000  38.375000 ;
      RECT  7.085000  38.305000 13.499000  38.375000 ;
      RECT  7.085000  38.375000 13.429000  38.445000 ;
      RECT  7.085000  38.375000 13.429000  38.445000 ;
      RECT  7.085000  38.445000 13.359000  38.515000 ;
      RECT  7.085000  38.445000 13.359000  38.515000 ;
      RECT  7.085000  38.515000 13.289000  38.585000 ;
      RECT  7.085000  38.515000 13.289000  38.585000 ;
      RECT  7.085000  38.585000 13.219000  38.655000 ;
      RECT  7.085000  38.585000 13.219000  38.655000 ;
      RECT  7.085000  38.655000 13.149000  38.725000 ;
      RECT  7.085000  38.655000 13.149000  38.725000 ;
      RECT  7.085000  38.725000 13.079000  38.795000 ;
      RECT  7.085000  38.725000 13.079000  38.795000 ;
      RECT  7.085000  38.795000 13.009000  38.865000 ;
      RECT  7.085000  38.795000 13.009000  38.865000 ;
      RECT  7.085000  38.865000 12.939000  38.935000 ;
      RECT  7.085000  38.865000 12.939000  38.935000 ;
      RECT  7.085000  38.935000 12.869000  39.005000 ;
      RECT  7.085000  38.935000 12.869000  39.005000 ;
      RECT  7.085000  39.005000 12.839000  39.035000 ;
      RECT  7.085000  39.005000 12.839000  39.035000 ;
      RECT  7.085000  39.036000 12.769000  39.105000 ;
      RECT  7.085000  39.036000 12.769000  39.105000 ;
      RECT  7.086000   9.255000 13.690000   9.310000 ;
      RECT  7.086000   9.255000 13.690000   9.310000 ;
      RECT  7.091000   1.675000 12.475000   1.745000 ;
      RECT  7.091000   1.675000 12.475000   1.745000 ;
      RECT  7.161000   1.745000 12.475000   1.815000 ;
      RECT  7.161000   1.745000 12.475000   1.815000 ;
      RECT  7.231000   1.815000 12.475000   1.885000 ;
      RECT  7.231000   1.815000 12.475000   1.885000 ;
      RECT  7.301000   1.885000 12.475000   1.955000 ;
      RECT  7.301000   1.885000 12.475000   1.955000 ;
      RECT  7.371000   1.955000 12.475000   2.025000 ;
      RECT  7.371000   1.955000 12.475000   2.025000 ;
      RECT  7.441000   2.025000 12.475000   2.095000 ;
      RECT  7.441000   2.025000 12.475000   2.095000 ;
      RECT  7.511000   2.095000 12.475000   2.165000 ;
      RECT  7.511000   2.095000 12.475000   2.165000 ;
      RECT  7.581000   2.165000 12.475000   2.235000 ;
      RECT  7.581000   2.165000 12.475000   2.235000 ;
      RECT  7.651000   2.235000 12.475000   2.305000 ;
      RECT  7.651000   2.235000 12.475000   2.305000 ;
      RECT  7.715000  56.628000 14.210000  57.837000 ;
      RECT  7.715000  57.837000 14.055000  57.992000 ;
      RECT  7.715000  57.992000 14.055000  58.450000 ;
      RECT  7.715000  58.450000 76.775000  73.557000 ;
      RECT  7.715000  73.557000 76.775000  74.047000 ;
      RECT  7.721000   2.305000 12.475000   2.375000 ;
      RECT  7.721000   2.305000 12.475000   2.375000 ;
      RECT  7.791000   2.375000 12.475000   2.445000 ;
      RECT  7.791000   2.375000 12.475000   2.445000 ;
      RECT  7.855000  56.686000 14.070000  57.779000 ;
      RECT  7.855000  57.779000 13.915000  73.499000 ;
      RECT  7.855000  57.779000 13.915000  73.499000 ;
      RECT  7.855000  57.779000 13.915000  73.499000 ;
      RECT  7.855000  57.779000 13.915000  73.499000 ;
      RECT  7.855000  57.779000 13.915000  73.499000 ;
      RECT  7.855000  57.779000 13.915000  73.499000 ;
      RECT  7.855000  57.779000 13.999000  57.850000 ;
      RECT  7.855000  57.779000 13.999000  57.850000 ;
      RECT  7.855000  57.850000 13.929000  57.920000 ;
      RECT  7.855000  57.850000 13.929000  57.920000 ;
      RECT  7.855000  57.920000 13.914000  57.935000 ;
      RECT  7.855000  57.920000 13.914000  57.935000 ;
      RECT  7.855000  57.934000 13.915000  58.590000 ;
      RECT  7.855000  58.590000 76.635000  73.499000 ;
      RECT  7.861000   2.445000 12.475000   2.515000 ;
      RECT  7.861000   2.445000 12.475000   2.515000 ;
      RECT  7.886000  56.655000 14.070000  56.685000 ;
      RECT  7.886000  56.655000 14.070000  56.685000 ;
      RECT  7.926000  73.499000 76.635000  73.570000 ;
      RECT  7.926000  73.499000 76.635000  73.570000 ;
      RECT  7.931000   2.515000 12.475000   2.585000 ;
      RECT  7.931000   2.515000 12.475000   2.585000 ;
      RECT  7.956000  56.585000 14.070000  56.655000 ;
      RECT  7.956000  56.585000 14.070000  56.655000 ;
      RECT  7.996000  73.570000 76.635000  73.640000 ;
      RECT  7.996000  73.570000 76.635000  73.640000 ;
      RECT  8.001000   2.585000 12.475000   2.655000 ;
      RECT  8.001000   2.585000 12.475000   2.655000 ;
      RECT  8.026000  56.515000 14.070000  56.585000 ;
      RECT  8.026000  56.515000 14.070000  56.585000 ;
      RECT  8.066000  73.640000 76.635000  73.710000 ;
      RECT  8.066000  73.640000 76.635000  73.710000 ;
      RECT  8.071000   2.655000 12.475000   2.725000 ;
      RECT  8.071000   2.655000 12.475000   2.725000 ;
      RECT  8.096000  56.445000 14.070000  56.515000 ;
      RECT  8.096000  56.445000 14.070000  56.515000 ;
      RECT  8.136000  73.710000 76.635000  73.780000 ;
      RECT  8.136000  73.710000 76.635000  73.780000 ;
      RECT  8.141000   2.725000 12.475000   2.795000 ;
      RECT  8.141000   2.725000 12.475000   2.795000 ;
      RECT  8.166000  56.375000 14.070000  56.445000 ;
      RECT  8.166000  56.375000 14.070000  56.445000 ;
      RECT  8.205000  74.047000 76.775000  74.622000 ;
      RECT  8.205000  74.622000 76.775000  75.027000 ;
      RECT  8.206000  73.780000 76.635000  73.850000 ;
      RECT  8.206000  73.780000 76.635000  73.850000 ;
      RECT  8.211000   2.795000 12.475000   2.865000 ;
      RECT  8.211000   2.795000 12.475000   2.865000 ;
      RECT  8.236000  56.305000 14.070000  56.375000 ;
      RECT  8.236000  56.305000 14.070000  56.375000 ;
      RECT  8.276000  73.850000 76.635000  73.920000 ;
      RECT  8.276000  73.850000 76.635000  73.920000 ;
      RECT  8.281000   2.865000 12.475000   2.935000 ;
      RECT  8.281000   2.865000 12.475000   2.935000 ;
      RECT  8.306000  56.235000 14.070000  56.305000 ;
      RECT  8.306000  56.235000 14.070000  56.305000 ;
      RECT  8.345000  73.989000 76.635000  74.564000 ;
      RECT  8.346000  73.920000 76.635000  73.990000 ;
      RECT  8.346000  73.920000 76.635000  73.990000 ;
      RECT  8.351000   2.935000 12.475000   3.005000 ;
      RECT  8.351000   2.935000 12.475000   3.005000 ;
      RECT  8.375000  54.128000 14.210000  55.968000 ;
      RECT  8.375000  55.968000 14.210000  56.628000 ;
      RECT  8.376000  56.165000 14.070000  56.235000 ;
      RECT  8.376000  56.165000 14.070000  56.235000 ;
      RECT  8.416000  74.564000 76.635000  74.635000 ;
      RECT  8.416000  74.564000 76.635000  74.635000 ;
      RECT  8.421000   3.005000 12.475000   3.075000 ;
      RECT  8.421000   3.005000 12.475000   3.075000 ;
      RECT  8.446000  56.095000 14.070000  56.165000 ;
      RECT  8.446000  56.095000 14.070000  56.165000 ;
      RECT  8.486000  74.635000 76.635000  74.705000 ;
      RECT  8.486000  74.635000 76.635000  74.705000 ;
      RECT  8.491000   3.075000 12.475000   3.145000 ;
      RECT  8.491000   3.075000 12.475000   3.145000 ;
      RECT  8.515000  54.186000 14.070000  56.026000 ;
      RECT  8.515000  56.026000 14.070000  56.095000 ;
      RECT  8.515000  56.026000 14.070000  56.095000 ;
      RECT  8.526000  54.175000 14.070000  54.185000 ;
      RECT  8.526000  54.175000 14.070000  54.185000 ;
      RECT  8.556000  74.705000 76.635000  74.775000 ;
      RECT  8.556000  74.705000 76.635000  74.775000 ;
      RECT  8.561000   3.145000 12.475000   3.215000 ;
      RECT  8.561000   3.145000 12.475000   3.215000 ;
      RECT  8.595000  44.243000 11.110000  47.443000 ;
      RECT  8.595000  47.443000 11.882000  48.215000 ;
      RECT  8.595000  48.215000 14.210000  48.743000 ;
      RECT  8.595000  48.743000 14.210000  53.908000 ;
      RECT  8.595000  53.908000 14.210000  54.128000 ;
      RECT  8.596000  54.105000 14.070000  54.175000 ;
      RECT  8.596000  54.105000 14.070000  54.175000 ;
      RECT  8.610000  75.027000 76.775000  77.137000 ;
      RECT  8.610000  77.137000 76.775000  77.227000 ;
      RECT  8.626000  74.775000 76.635000  74.845000 ;
      RECT  8.626000  74.775000 76.635000  74.845000 ;
      RECT  8.631000   3.215000 12.475000   3.285000 ;
      RECT  8.631000   3.215000 12.475000   3.285000 ;
      RECT  8.666000  54.035000 14.070000  54.105000 ;
      RECT  8.666000  54.035000 14.070000  54.105000 ;
      RECT  8.696000  74.845000 76.635000  74.915000 ;
      RECT  8.696000  74.845000 76.635000  74.915000 ;
      RECT  8.700000  77.227000 76.775000  77.685000 ;
      RECT  8.701000   3.285000 12.475000   3.355000 ;
      RECT  8.701000   3.285000 12.475000   3.355000 ;
      RECT  8.735000  44.301000 10.970000  45.266000 ;
      RECT  8.735000  45.335000  8.804000  45.405000 ;
      RECT  8.735000  45.335000  8.804000  45.405000 ;
      RECT  8.735000  45.405000  8.874000  45.475000 ;
      RECT  8.735000  45.405000  8.874000  45.475000 ;
      RECT  8.735000  45.475000  8.944000  45.545000 ;
      RECT  8.735000  45.475000  8.944000  45.545000 ;
      RECT  8.735000  45.545000  9.014000  45.615000 ;
      RECT  8.735000  45.545000  9.014000  45.615000 ;
      RECT  8.735000  45.615000  9.084000  45.685000 ;
      RECT  8.735000  45.615000  9.084000  45.685000 ;
      RECT  8.735000  45.685000  9.154000  45.755000 ;
      RECT  8.735000  45.685000  9.154000  45.755000 ;
      RECT  8.735000  45.755000  9.224000  45.825000 ;
      RECT  8.735000  45.755000  9.224000  45.825000 ;
      RECT  8.735000  45.825000  9.294000  45.895000 ;
      RECT  8.735000  45.825000  9.294000  45.895000 ;
      RECT  8.735000  45.895000  9.364000  45.965000 ;
      RECT  8.735000  45.895000  9.364000  45.965000 ;
      RECT  8.735000  45.965000  9.434000  46.035000 ;
      RECT  8.735000  45.965000  9.434000  46.035000 ;
      RECT  8.735000  46.035000  9.504000  46.105000 ;
      RECT  8.735000  46.035000  9.504000  46.105000 ;
      RECT  8.735000  46.105000  9.574000  46.175000 ;
      RECT  8.735000  46.105000  9.574000  46.175000 ;
      RECT  8.735000  46.175000  9.644000  46.245000 ;
      RECT  8.735000  46.175000  9.644000  46.245000 ;
      RECT  8.735000  46.245000  9.714000  46.315000 ;
      RECT  8.735000  46.245000  9.714000  46.315000 ;
      RECT  8.735000  46.315000  9.784000  46.385000 ;
      RECT  8.735000  46.315000  9.784000  46.385000 ;
      RECT  8.735000  46.385000  9.854000  46.455000 ;
      RECT  8.735000  46.385000  9.854000  46.455000 ;
      RECT  8.735000  46.455000  9.924000  46.525000 ;
      RECT  8.735000  46.455000  9.924000  46.525000 ;
      RECT  8.735000  46.525000  9.994000  46.595000 ;
      RECT  8.735000  46.525000  9.994000  46.595000 ;
      RECT  8.735000  46.595000 10.064000  46.665000 ;
      RECT  8.735000  46.595000 10.064000  46.665000 ;
      RECT  8.735000  46.665000 10.134000  46.735000 ;
      RECT  8.735000  46.665000 10.134000  46.735000 ;
      RECT  8.735000  46.735000 10.204000  46.805000 ;
      RECT  8.735000  46.735000 10.204000  46.805000 ;
      RECT  8.735000  46.805000 10.274000  46.875000 ;
      RECT  8.735000  46.805000 10.274000  46.875000 ;
      RECT  8.735000  46.875000 10.344000  46.945000 ;
      RECT  8.735000  46.875000 10.344000  46.945000 ;
      RECT  8.735000  46.945000 10.414000  47.015000 ;
      RECT  8.735000  46.945000 10.414000  47.015000 ;
      RECT  8.735000  47.015000 10.484000  47.085000 ;
      RECT  8.735000  47.015000 10.484000  47.085000 ;
      RECT  8.735000  47.085000 10.554000  47.155000 ;
      RECT  8.735000  47.085000 10.554000  47.155000 ;
      RECT  8.735000  47.155000 10.624000  47.225000 ;
      RECT  8.735000  47.155000 10.624000  47.225000 ;
      RECT  8.735000  47.225000 10.694000  47.295000 ;
      RECT  8.735000  47.225000 10.694000  47.295000 ;
      RECT  8.735000  47.295000 10.764000  47.365000 ;
      RECT  8.735000  47.295000 10.764000  47.365000 ;
      RECT  8.735000  47.365000 10.834000  47.435000 ;
      RECT  8.735000  47.365000 10.834000  47.435000 ;
      RECT  8.735000  47.435000 10.904000  47.500000 ;
      RECT  8.735000  47.435000 10.904000  47.500000 ;
      RECT  8.735000  47.501000 10.970000  47.570000 ;
      RECT  8.735000  47.501000 10.970000  47.570000 ;
      RECT  8.735000  47.570000 11.039000  47.640000 ;
      RECT  8.735000  47.570000 11.039000  47.640000 ;
      RECT  8.735000  47.640000 11.109000  47.710000 ;
      RECT  8.735000  47.640000 11.109000  47.710000 ;
      RECT  8.735000  47.710000 11.179000  47.780000 ;
      RECT  8.735000  47.710000 11.179000  47.780000 ;
      RECT  8.735000  47.780000 11.249000  47.850000 ;
      RECT  8.735000  47.780000 11.249000  47.850000 ;
      RECT  8.735000  47.850000 11.319000  47.920000 ;
      RECT  8.735000  47.850000 11.319000  47.920000 ;
      RECT  8.735000  47.920000 11.389000  47.990000 ;
      RECT  8.735000  47.920000 11.389000  47.990000 ;
      RECT  8.735000  47.990000 11.459000  48.060000 ;
      RECT  8.735000  47.990000 11.459000  48.060000 ;
      RECT  8.735000  48.060000 11.529000  48.130000 ;
      RECT  8.735000  48.060000 11.529000  48.130000 ;
      RECT  8.735000  48.130000 11.599000  48.200000 ;
      RECT  8.735000  48.130000 11.599000  48.200000 ;
      RECT  8.735000  48.200000 11.669000  48.270000 ;
      RECT  8.735000  48.200000 11.669000  48.270000 ;
      RECT  8.735000  48.270000 11.739000  48.340000 ;
      RECT  8.735000  48.270000 11.739000  48.340000 ;
      RECT  8.735000  48.340000 11.809000  48.355000 ;
      RECT  8.735000  48.340000 11.809000  48.355000 ;
      RECT  8.735000  48.355000 13.624000  48.425000 ;
      RECT  8.735000  48.355000 13.624000  48.425000 ;
      RECT  8.735000  48.425000 13.694000  48.495000 ;
      RECT  8.735000  48.425000 13.694000  48.495000 ;
      RECT  8.735000  48.495000 13.764000  48.565000 ;
      RECT  8.735000  48.495000 13.764000  48.565000 ;
      RECT  8.735000  48.565000 13.834000  48.635000 ;
      RECT  8.735000  48.565000 13.834000  48.635000 ;
      RECT  8.735000  48.635000 13.904000  48.705000 ;
      RECT  8.735000  48.635000 13.904000  48.705000 ;
      RECT  8.735000  48.705000 13.974000  48.775000 ;
      RECT  8.735000  48.705000 13.974000  48.775000 ;
      RECT  8.735000  48.775000 14.044000  48.800000 ;
      RECT  8.735000  48.775000 14.044000  48.800000 ;
      RECT  8.735000  48.801000 14.070000  53.966000 ;
      RECT  8.735000  48.801000 14.070000  56.026000 ;
      RECT  8.735000  48.801000 14.070000  56.686000 ;
      RECT  8.735000  48.801000 14.070000  56.686000 ;
      RECT  8.735000  48.801000 14.070000  56.686000 ;
      RECT  8.735000  48.801000 14.070000  56.686000 ;
      RECT  8.735000  53.966000 14.070000  54.035000 ;
      RECT  8.735000  53.966000 14.070000  54.035000 ;
      RECT  8.750000  74.969000 76.635000  77.079000 ;
      RECT  8.751000  74.915000 76.635000  74.970000 ;
      RECT  8.751000  74.915000 76.635000  74.970000 ;
      RECT  8.756000  44.280000 10.970000  44.300000 ;
      RECT  8.771000   3.355000 12.475000   3.425000 ;
      RECT  8.771000   3.355000 12.475000   3.425000 ;
      RECT  8.796000  77.079000 76.635000  77.125000 ;
      RECT  8.796000  77.079000 76.635000  77.125000 ;
      RECT  8.826000  44.210000 10.970000  44.280000 ;
      RECT  8.840000  74.969000 76.635000  96.079000 ;
      RECT  8.840000  74.969000 76.635000  96.079000 ;
      RECT  8.841000   3.425000 12.475000   3.495000 ;
      RECT  8.841000   3.425000 12.475000   3.495000 ;
      RECT  8.841000  77.125000 76.635000  77.170000 ;
      RECT  8.841000  77.125000 76.635000  77.170000 ;
      RECT  8.845000   3.697000 12.615000   5.408000 ;
      RECT  8.845000   5.408000 13.830000   6.623000 ;
      RECT  8.845000   6.623000 13.830000   6.920000 ;
      RECT  8.896000  44.140000 10.970000  44.210000 ;
      RECT  8.911000   3.495000 12.475000   3.565000 ;
      RECT  8.911000   3.495000 12.475000   3.565000 ;
      RECT  8.966000  44.070000 10.970000  44.140000 ;
      RECT  8.981000   3.565000 12.475000   3.635000 ;
      RECT  8.981000   3.565000 12.475000   3.635000 ;
      RECT  8.985000   1.324000 12.475000   5.466000 ;
      RECT  8.985000   1.324000 12.475000   5.466000 ;
      RECT  8.985000   1.324000 12.475000   5.466000 ;
      RECT  8.985000   1.324000 12.475000   5.466000 ;
      RECT  8.985000   5.466000 12.475000   5.535000 ;
      RECT  8.985000   5.466000 12.475000   5.535000 ;
      RECT  8.985000   5.535000 12.544000   5.605000 ;
      RECT  8.985000   5.535000 12.544000   5.605000 ;
      RECT  8.985000   5.605000 12.614000   5.675000 ;
      RECT  8.985000   5.605000 12.614000   5.675000 ;
      RECT  8.985000   5.675000 12.684000   5.745000 ;
      RECT  8.985000   5.675000 12.684000   5.745000 ;
      RECT  8.985000   5.745000 12.754000   5.815000 ;
      RECT  8.985000   5.745000 12.754000   5.815000 ;
      RECT  8.985000   5.815000 12.824000   5.885000 ;
      RECT  8.985000   5.815000 12.824000   5.885000 ;
      RECT  8.985000   5.885000 12.894000   5.955000 ;
      RECT  8.985000   5.885000 12.894000   5.955000 ;
      RECT  8.985000   5.955000 12.964000   6.025000 ;
      RECT  8.985000   5.955000 12.964000   6.025000 ;
      RECT  8.985000   6.025000 13.034000   6.095000 ;
      RECT  8.985000   6.025000 13.034000   6.095000 ;
      RECT  8.985000   6.095000 13.104000   6.165000 ;
      RECT  8.985000   6.095000 13.104000   6.165000 ;
      RECT  8.985000   6.165000 13.174000   6.235000 ;
      RECT  8.985000   6.165000 13.174000   6.235000 ;
      RECT  8.985000   6.235000 13.244000   6.305000 ;
      RECT  8.985000   6.235000 13.244000   6.305000 ;
      RECT  8.985000   6.305000 13.314000   6.375000 ;
      RECT  8.985000   6.305000 13.314000   6.375000 ;
      RECT  8.985000   6.375000 13.384000   6.445000 ;
      RECT  8.985000   6.375000 13.384000   6.445000 ;
      RECT  8.985000   6.445000 13.454000   6.515000 ;
      RECT  8.985000   6.445000 13.454000   6.515000 ;
      RECT  8.985000   6.515000 13.524000   6.585000 ;
      RECT  8.985000   6.515000 13.524000   6.585000 ;
      RECT  8.985000   6.585000 13.594000   6.655000 ;
      RECT  8.985000   6.585000 13.594000   6.655000 ;
      RECT  8.985000   6.655000 13.664000   6.680000 ;
      RECT  8.985000   6.655000 13.664000   6.680000 ;
      RECT  8.985000   6.681000 13.690000   7.060000 ;
      RECT  8.986000   3.635000 12.475000   3.640000 ;
      RECT  8.986000   3.635000 12.475000   3.640000 ;
      RECT  9.036000  44.000000 10.970000  44.070000 ;
      RECT  9.061000  43.777000 11.110000  44.243000 ;
      RECT  9.106000  43.930000 10.970000  44.000000 ;
      RECT  9.176000  43.860000 10.970000  43.930000 ;
      RECT  9.246000  43.790000 10.970000  43.860000 ;
      RECT  9.317000  43.719000 10.970000  43.790000 ;
      RECT  9.376000  43.660000 10.969000  43.720000 ;
      RECT  9.446000  43.590000 11.029000  43.660000 ;
      RECT  9.516000  43.520000 11.099000  43.590000 ;
      RECT  9.586000  43.450000 11.169000  43.520000 ;
      RECT  9.656000  43.380000 11.239000  43.450000 ;
      RECT  9.726000  43.310000 11.309000  43.380000 ;
      RECT  9.796000  43.240000 11.379000  43.310000 ;
      RECT  9.866000  43.170000 11.449000  43.240000 ;
      RECT  9.936000  43.100000 11.519000  43.170000 ;
      RECT 10.006000  43.030000 11.589000  43.100000 ;
      RECT 10.076000  42.960000 11.659000  43.030000 ;
      RECT 10.146000  42.890000 11.729000  42.960000 ;
      RECT 10.216000  42.820000 11.799000  42.890000 ;
      RECT 10.286000  42.750000 11.869000  42.820000 ;
      RECT 10.356000  42.680000 11.939000  42.750000 ;
      RECT 10.426000  42.610000 12.009000  42.680000 ;
      RECT 10.496000  42.540000 12.079000  42.610000 ;
      RECT 10.566000  42.470000 12.149000  42.540000 ;
      RECT 10.636000  42.400000 12.219000  42.470000 ;
      RECT 10.706000  42.330000 12.289000  42.400000 ;
      RECT 10.776000  42.260000 12.359000  42.330000 ;
      RECT 10.846000  42.190000 12.429000  42.260000 ;
      RECT 10.916000  42.120000 12.499000  42.190000 ;
      RECT 10.986000  42.050000 12.569000  42.120000 ;
      RECT 11.056000  41.980000 12.639000  42.050000 ;
      RECT 11.126000  41.910000 12.709000  41.980000 ;
      RECT 11.196000  41.840000 12.779000  41.910000 ;
      RECT 11.266000  41.770000 12.849000  41.840000 ;
      RECT 11.336000  41.700000 12.919000  41.770000 ;
      RECT 11.406000  41.630000 12.989000  41.700000 ;
      RECT 11.476000  41.560000 13.059000  41.630000 ;
      RECT 11.546000  41.490000 13.129000  41.560000 ;
      RECT 11.616000  41.420000 13.199000  41.490000 ;
      RECT 11.650000  44.003000 29.985000  47.217000 ;
      RECT 11.650000  47.217000 29.985000  47.675000 ;
      RECT 11.687000  41.349000 13.269000  41.420000 ;
      RECT 11.741000  41.295000 13.340000  41.350000 ;
      RECT 11.790000  44.061000 29.845000  47.159000 ;
      RECT 11.811000  41.225000 13.340000  41.295000 ;
      RECT 11.851000  44.000000 29.845000  44.060000 ;
      RECT 11.851000  44.000000 29.845000  44.060000 ;
      RECT 11.861000  47.159000 29.845000  47.230000 ;
      RECT 11.861000  47.159000 29.845000  47.230000 ;
      RECT 11.881000  41.155000 13.340000  41.225000 ;
      RECT 11.921000  43.930000 29.845000  44.000000 ;
      RECT 11.921000  43.930000 29.845000  44.000000 ;
      RECT 11.931000  47.230000 29.845000  47.300000 ;
      RECT 11.931000  47.230000 29.845000  47.300000 ;
      RECT 11.951000  41.085000 13.340000  41.155000 ;
      RECT 11.991000  43.860000 29.845000  43.930000 ;
      RECT 11.991000  43.860000 29.845000  43.930000 ;
      RECT 12.001000  47.300000 29.845000  47.370000 ;
      RECT 12.001000  47.300000 29.845000  47.370000 ;
      RECT 12.021000  41.015000 13.340000  41.085000 ;
      RECT 12.061000  43.790000 29.845000  43.860000 ;
      RECT 12.061000  43.790000 29.845000  43.860000 ;
      RECT 12.071000  47.370000 29.845000  47.440000 ;
      RECT 12.071000  47.370000 29.845000  47.440000 ;
      RECT 12.091000  40.945000 13.340000  41.015000 ;
      RECT 12.131000  43.720000 29.845000  43.790000 ;
      RECT 12.131000  43.720000 29.845000  43.790000 ;
      RECT 12.141000  47.440000 29.845000  47.510000 ;
      RECT 12.141000  47.440000 29.845000  47.510000 ;
      RECT 12.161000  40.875000 13.340000  40.945000 ;
      RECT 12.166000  47.510000 29.845000  47.535000 ;
      RECT 12.166000  47.510000 29.845000  47.535000 ;
      RECT 12.201000  43.650000 29.845000  43.720000 ;
      RECT 12.201000  43.650000 29.845000  43.720000 ;
      RECT 12.231000  40.805000 13.340000  40.875000 ;
      RECT 12.271000  43.580000 29.845000  43.650000 ;
      RECT 12.271000  43.580000 29.845000  43.650000 ;
      RECT 12.301000  40.735000 13.340000  40.805000 ;
      RECT 12.341000  43.510000 29.845000  43.580000 ;
      RECT 12.341000  43.510000 29.845000  43.580000 ;
      RECT 12.371000  40.665000 13.340000  40.735000 ;
      RECT 12.411000  43.440000 29.845000  43.510000 ;
      RECT 12.411000  43.440000 29.845000  43.510000 ;
      RECT 12.441000  40.595000 13.340000  40.665000 ;
      RECT 12.466000  40.372000 13.480000  41.407000 ;
      RECT 12.481000  43.370000 29.845000  43.440000 ;
      RECT 12.481000  43.370000 29.845000  43.440000 ;
      RECT 12.511000  40.525000 13.340000  40.595000 ;
      RECT 12.551000  43.300000 29.845000  43.370000 ;
      RECT 12.551000  43.300000 29.845000  43.370000 ;
      RECT 12.581000  40.455000 13.340000  40.525000 ;
      RECT 12.621000  43.230000 29.845000  43.300000 ;
      RECT 12.621000  43.230000 29.845000  43.300000 ;
      RECT 12.651000  40.385000 13.340000  40.455000 ;
      RECT 12.691000  43.160000 29.845000  43.230000 ;
      RECT 12.691000  43.160000 29.845000  43.230000 ;
      RECT 12.722000  40.314000 13.340000  40.385000 ;
      RECT 12.746000  40.290000 13.339000  40.315000 ;
      RECT 12.761000  43.090000 29.845000  43.160000 ;
      RECT 12.761000  43.090000 29.845000  43.160000 ;
      RECT 12.816000  40.220000 13.364000  40.290000 ;
      RECT 12.831000  43.020000 29.845000  43.090000 ;
      RECT 12.831000  43.020000 29.845000  43.090000 ;
      RECT 12.886000  40.150000 13.434000  40.220000 ;
      RECT 12.901000  42.950000 29.845000  43.020000 ;
      RECT 12.901000  42.950000 29.845000  43.020000 ;
      RECT 12.956000  40.080000 13.504000  40.150000 ;
      RECT 12.971000  42.880000 29.845000  42.950000 ;
      RECT 12.971000  42.880000 29.845000  42.950000 ;
      RECT 13.026000  40.010000 13.574000  40.080000 ;
      RECT 13.041000  42.810000 29.845000  42.880000 ;
      RECT 13.041000  42.810000 29.845000  42.880000 ;
      RECT 13.096000  39.940000 13.644000  40.010000 ;
      RECT 13.111000  42.740000 29.845000  42.810000 ;
      RECT 13.111000  42.740000 29.845000  42.810000 ;
      RECT 13.155000   0.000000 16.170000   2.378000 ;
      RECT 13.155000   2.378000 16.955000   3.163000 ;
      RECT 13.155000   3.163000 16.955000   5.182000 ;
      RECT 13.155000   5.182000 16.955000   6.397000 ;
      RECT 13.166000  39.870000 13.714000  39.940000 ;
      RECT 13.181000  42.670000 29.845000  42.740000 ;
      RECT 13.181000  42.670000 29.845000  42.740000 ;
      RECT 13.236000  39.800000 13.784000  39.870000 ;
      RECT 13.251000  42.600000 29.845000  42.670000 ;
      RECT 13.251000  42.600000 29.845000  42.670000 ;
      RECT 13.295000   0.000000 13.594000   0.070000 ;
      RECT 13.295000   0.000000 13.594000   0.070000 ;
      RECT 13.295000   0.070000 13.664000   0.140000 ;
      RECT 13.295000   0.070000 13.664000   0.140000 ;
      RECT 13.295000   0.140000 13.734000   0.210000 ;
      RECT 13.295000   0.140000 13.734000   0.210000 ;
      RECT 13.295000   0.210000 13.804000   0.280000 ;
      RECT 13.295000   0.210000 13.804000   0.280000 ;
      RECT 13.295000   0.280000 13.874000   0.350000 ;
      RECT 13.295000   0.280000 13.874000   0.350000 ;
      RECT 13.295000   0.350000 13.944000   0.420000 ;
      RECT 13.295000   0.350000 13.944000   0.420000 ;
      RECT 13.295000   0.420000 14.014000   0.490000 ;
      RECT 13.295000   0.420000 14.014000   0.490000 ;
      RECT 13.295000   0.490000 14.084000   0.560000 ;
      RECT 13.295000   0.490000 14.084000   0.560000 ;
      RECT 13.295000   0.560000 14.154000   0.630000 ;
      RECT 13.295000   0.560000 14.154000   0.630000 ;
      RECT 13.295000   0.630000 14.224000   0.700000 ;
      RECT 13.295000   0.630000 14.224000   0.700000 ;
      RECT 13.295000   0.700000 14.294000   0.770000 ;
      RECT 13.295000   0.700000 14.294000   0.770000 ;
      RECT 13.295000   0.770000 14.364000   0.840000 ;
      RECT 13.295000   0.770000 14.364000   0.840000 ;
      RECT 13.295000   0.840000 14.434000   0.910000 ;
      RECT 13.295000   0.840000 14.434000   0.910000 ;
      RECT 13.295000   0.910000 14.504000   0.980000 ;
      RECT 13.295000   0.910000 14.504000   0.980000 ;
      RECT 13.295000   0.980000 14.574000   1.050000 ;
      RECT 13.295000   0.980000 14.574000   1.050000 ;
      RECT 13.295000   1.050000 14.644000   1.120000 ;
      RECT 13.295000   1.050000 14.644000   1.120000 ;
      RECT 13.295000   1.120000 14.714000   1.190000 ;
      RECT 13.295000   1.120000 14.714000   1.190000 ;
      RECT 13.295000   1.190000 14.784000   1.260000 ;
      RECT 13.295000   1.190000 14.784000   1.260000 ;
      RECT 13.295000   1.260000 14.854000   1.330000 ;
      RECT 13.295000   1.260000 14.854000   1.330000 ;
      RECT 13.295000   1.330000 14.924000   1.400000 ;
      RECT 13.295000   1.330000 14.924000   1.400000 ;
      RECT 13.295000   1.400000 14.994000   1.470000 ;
      RECT 13.295000   1.400000 14.994000   1.470000 ;
      RECT 13.295000   1.470000 15.064000   1.540000 ;
      RECT 13.295000   1.470000 15.064000   1.540000 ;
      RECT 13.295000   1.540000 15.134000   1.610000 ;
      RECT 13.295000   1.540000 15.134000   1.610000 ;
      RECT 13.295000   1.610000 15.204000   1.680000 ;
      RECT 13.295000   1.610000 15.204000   1.680000 ;
      RECT 13.295000   1.680000 15.274000   1.750000 ;
      RECT 13.295000   1.680000 15.274000   1.750000 ;
      RECT 13.295000   1.750000 15.344000   1.820000 ;
      RECT 13.295000   1.750000 15.344000   1.820000 ;
      RECT 13.295000   1.820000 15.414000   1.890000 ;
      RECT 13.295000   1.820000 15.414000   1.890000 ;
      RECT 13.295000   1.890000 15.484000   1.960000 ;
      RECT 13.295000   1.890000 15.484000   1.960000 ;
      RECT 13.295000   1.960000 15.554000   2.030000 ;
      RECT 13.295000   1.960000 15.554000   2.030000 ;
      RECT 13.295000   2.030000 15.624000   2.100000 ;
      RECT 13.295000   2.030000 15.624000   2.100000 ;
      RECT 13.295000   2.100000 15.694000   2.170000 ;
      RECT 13.295000   2.100000 15.694000   2.170000 ;
      RECT 13.295000   2.170000 15.764000   2.240000 ;
      RECT 13.295000   2.170000 15.764000   2.240000 ;
      RECT 13.295000   2.240000 15.834000   2.310000 ;
      RECT 13.295000   2.240000 15.834000   2.310000 ;
      RECT 13.295000   2.310000 15.904000   2.380000 ;
      RECT 13.295000   2.310000 15.904000   2.380000 ;
      RECT 13.295000   2.380000 15.974000   2.435000 ;
      RECT 13.295000   2.380000 15.974000   2.435000 ;
      RECT 13.295000   2.436000 16.030000   2.505000 ;
      RECT 13.295000   2.436000 16.030000   2.505000 ;
      RECT 13.295000   2.505000 16.099000   2.575000 ;
      RECT 13.295000   2.505000 16.099000   2.575000 ;
      RECT 13.295000   2.575000 16.169000   2.645000 ;
      RECT 13.295000   2.575000 16.169000   2.645000 ;
      RECT 13.295000   2.645000 16.239000   2.715000 ;
      RECT 13.295000   2.645000 16.239000   2.715000 ;
      RECT 13.295000   2.715000 16.309000   2.785000 ;
      RECT 13.295000   2.715000 16.309000   2.785000 ;
      RECT 13.295000   2.785000 16.379000   2.855000 ;
      RECT 13.295000   2.785000 16.379000   2.855000 ;
      RECT 13.295000   2.855000 16.449000   2.925000 ;
      RECT 13.295000   2.855000 16.449000   2.925000 ;
      RECT 13.295000   2.925000 16.519000   2.995000 ;
      RECT 13.295000   2.925000 16.519000   2.995000 ;
      RECT 13.295000   2.995000 16.589000   3.065000 ;
      RECT 13.295000   2.995000 16.589000   3.065000 ;
      RECT 13.295000   3.065000 16.659000   3.135000 ;
      RECT 13.295000   3.065000 16.659000   3.135000 ;
      RECT 13.295000   3.135000 16.729000   3.205000 ;
      RECT 13.295000   3.135000 16.729000   3.205000 ;
      RECT 13.295000   3.205000 16.799000   3.220000 ;
      RECT 13.295000   3.205000 16.799000   3.220000 ;
      RECT 13.295000   3.221000 16.815000   5.124000 ;
      RECT 13.306000  39.730000 13.854000  39.800000 ;
      RECT 13.318000  39.520000 13.480000  40.372000 ;
      RECT 13.321000  42.530000 29.845000  42.600000 ;
      RECT 13.321000  42.530000 29.845000  42.600000 ;
      RECT 13.366000   5.124000 16.815000   5.195000 ;
      RECT 13.366000   5.124000 16.815000   5.195000 ;
      RECT 13.376000  39.660000 13.924000  39.730000 ;
      RECT 13.391000  42.460000 29.845000  42.530000 ;
      RECT 13.391000  42.460000 29.845000  42.530000 ;
      RECT 13.436000   5.195000 16.815000   5.265000 ;
      RECT 13.436000   5.195000 16.815000   5.265000 ;
      RECT 13.446000  39.590000 13.994000  39.660000 ;
      RECT 13.461000  42.390000 29.845000  42.460000 ;
      RECT 13.461000  42.390000 29.845000  42.460000 ;
      RECT 13.506000   5.265000 16.815000   5.335000 ;
      RECT 13.506000   5.265000 16.815000   5.335000 ;
      RECT 13.516000  39.520000 14.064000  39.590000 ;
      RECT 13.531000  42.320000 29.845000  42.390000 ;
      RECT 13.531000  42.320000 29.845000  42.390000 ;
      RECT 13.576000   5.335000 16.815000   5.405000 ;
      RECT 13.576000   5.335000 16.815000   5.405000 ;
      RECT 13.586000  39.450000 14.134000  39.520000 ;
      RECT 13.601000  42.250000 29.845000  42.320000 ;
      RECT 13.601000  42.250000 29.845000  42.320000 ;
      RECT 13.646000   5.405000 16.815000   5.475000 ;
      RECT 13.646000   5.405000 16.815000   5.475000 ;
      RECT 13.656000  39.380000 14.204000  39.450000 ;
      RECT 13.671000  42.180000 29.845000  42.250000 ;
      RECT 13.671000  42.180000 29.845000  42.250000 ;
      RECT 13.691000  39.345000 15.194000  39.380000 ;
      RECT 13.716000   5.475000 16.815000   5.545000 ;
      RECT 13.716000   5.475000 16.815000   5.545000 ;
      RECT 13.741000  42.110000 29.845000  42.180000 ;
      RECT 13.741000  42.110000 29.845000  42.180000 ;
      RECT 13.761000  39.275000 15.229000  39.345000 ;
      RECT 13.786000   5.545000 16.815000   5.615000 ;
      RECT 13.786000   5.545000 16.815000   5.615000 ;
      RECT 13.811000  42.040000 29.845000  42.110000 ;
      RECT 13.811000  42.040000 29.845000  42.110000 ;
      RECT 13.831000  39.205000 15.299000  39.275000 ;
      RECT 13.856000   5.615000 16.815000   5.685000 ;
      RECT 13.856000   5.615000 16.815000   5.685000 ;
      RECT 13.881000  41.970000 29.845000  42.040000 ;
      RECT 13.881000  41.970000 29.845000  42.040000 ;
      RECT 13.901000  39.135000 15.369000  39.205000 ;
      RECT 13.908000  47.675000 29.985000  48.517000 ;
      RECT 13.926000   5.685000 16.815000   5.755000 ;
      RECT 13.926000   5.685000 16.815000   5.755000 ;
      RECT 13.951000  41.900000 29.845000  41.970000 ;
      RECT 13.951000  41.900000 29.845000  41.970000 ;
      RECT 13.971000  39.065000 15.439000  39.135000 ;
      RECT 13.996000   5.755000 16.815000   5.825000 ;
      RECT 13.996000   5.755000 16.815000   5.825000 ;
      RECT 14.020000  40.598000 29.985000  41.633000 ;
      RECT 14.020000  41.633000 29.985000  44.003000 ;
      RECT 14.021000  41.830000 29.845000  41.900000 ;
      RECT 14.021000  41.830000 29.845000  41.900000 ;
      RECT 14.036000  47.535000 29.845000  47.605000 ;
      RECT 14.036000  47.535000 29.845000  47.605000 ;
      RECT 14.041000  38.995000 15.509000  39.065000 ;
      RECT 14.066000   5.825000 16.815000   5.895000 ;
      RECT 14.066000   5.825000 16.815000   5.895000 ;
      RECT 14.091000  41.760000 29.845000  41.830000 ;
      RECT 14.091000  41.760000 29.845000  41.830000 ;
      RECT 14.106000  47.605000 29.845000  47.675000 ;
      RECT 14.106000  47.605000 29.845000  47.675000 ;
      RECT 14.111000  38.925000 15.579000  38.995000 ;
      RECT 14.136000   5.895000 16.815000   5.965000 ;
      RECT 14.136000   5.895000 16.815000   5.965000 ;
      RECT 14.160000  40.656000 29.845000  41.691000 ;
      RECT 14.160000  41.691000 29.845000  41.760000 ;
      RECT 14.160000  41.691000 29.845000  41.760000 ;
      RECT 14.176000  47.675000 29.845000  47.745000 ;
      RECT 14.176000  47.675000 29.845000  47.745000 ;
      RECT 14.181000  38.855000 15.649000  38.925000 ;
      RECT 14.196000  40.620000 29.845000  40.655000 ;
      RECT 14.196000  40.620000 29.845000  40.655000 ;
      RECT 14.206000   5.965000 16.815000   6.035000 ;
      RECT 14.206000   5.965000 16.815000   6.035000 ;
      RECT 14.246000  47.745000 29.845000  47.815000 ;
      RECT 14.246000  47.745000 29.845000  47.815000 ;
      RECT 14.251000  38.785000 15.719000  38.855000 ;
      RECT 14.266000  40.550000 29.845000  40.620000 ;
      RECT 14.266000  40.550000 29.845000  40.620000 ;
      RECT 14.276000   6.035000 16.815000   6.105000 ;
      RECT 14.276000   6.035000 16.815000   6.105000 ;
      RECT 14.316000  47.815000 29.845000  47.885000 ;
      RECT 14.316000  47.815000 29.845000  47.885000 ;
      RECT 14.321000  38.715000 15.789000  38.785000 ;
      RECT 14.336000  40.480000 29.845000  40.550000 ;
      RECT 14.336000  40.480000 29.845000  40.550000 ;
      RECT 14.346000   6.105000 16.815000   6.175000 ;
      RECT 14.346000   6.105000 16.815000   6.175000 ;
      RECT 14.370000   6.397000 16.955000   6.617000 ;
      RECT 14.370000   6.617000 16.470000   7.102000 ;
      RECT 14.370000   7.102000 16.470000  11.598000 ;
      RECT 14.370000  11.598000 16.565000  11.693000 ;
      RECT 14.370000  11.693000 16.565000  12.322000 ;
      RECT 14.370000  12.322000 16.470000  12.417000 ;
      RECT 14.370000  12.417000 16.470000  18.057000 ;
      RECT 14.370000  18.057000 16.470000  19.472000 ;
      RECT 14.386000  47.885000 29.845000  47.955000 ;
      RECT 14.386000  47.885000 29.845000  47.955000 ;
      RECT 14.391000  38.645000 15.859000  38.715000 ;
      RECT 14.406000  40.410000 29.845000  40.480000 ;
      RECT 14.406000  40.410000 29.845000  40.480000 ;
      RECT 14.416000   6.175000 16.815000   6.245000 ;
      RECT 14.416000   6.175000 16.815000   6.245000 ;
      RECT 14.456000  47.955000 29.845000  48.025000 ;
      RECT 14.456000  47.955000 29.845000  48.025000 ;
      RECT 14.461000  38.575000 15.929000  38.645000 ;
      RECT 14.476000  40.340000 29.845000  40.410000 ;
      RECT 14.476000  40.340000 29.845000  40.410000 ;
      RECT 14.486000   6.245000 16.815000   6.315000 ;
      RECT 14.486000   6.245000 16.815000   6.315000 ;
      RECT 14.510000   6.559000 16.744000   6.630000 ;
      RECT 14.510000   6.630000 16.674000   6.700000 ;
      RECT 14.510000   6.700000 16.604000   6.770000 ;
      RECT 14.510000   6.770000 16.534000   6.840000 ;
      RECT 14.510000   6.840000 16.464000   6.910000 ;
      RECT 14.510000   6.910000 16.394000   6.980000 ;
      RECT 14.510000   6.980000 16.329000   7.045000 ;
      RECT 14.510000   7.044000 16.330000  11.656000 ;
      RECT 14.510000  11.656000 16.330000  11.705000 ;
      RECT 14.510000  11.705000 16.379000  11.750000 ;
      RECT 14.510000  11.751000 16.425000  12.264000 ;
      RECT 14.510000  12.264000 16.379000  12.310000 ;
      RECT 14.510000  12.310000 16.334000  12.355000 ;
      RECT 14.510000  12.355000 16.329000  12.360000 ;
      RECT 14.510000  12.359000 16.330000  17.999000 ;
      RECT 14.511000   6.315000 16.815000   6.340000 ;
      RECT 14.511000   6.315000 16.815000   6.340000 ;
      RECT 14.526000  48.025000 29.845000  48.095000 ;
      RECT 14.526000  48.025000 29.845000  48.095000 ;
      RECT 14.531000  38.505000 15.999000  38.575000 ;
      RECT 14.546000  40.270000 29.845000  40.340000 ;
      RECT 14.546000  40.270000 29.845000  40.340000 ;
      RECT 14.558000  40.060000 29.985000  40.598000 ;
      RECT 14.581000   6.339000 16.815000   6.410000 ;
      RECT 14.581000   6.339000 16.815000   6.410000 ;
      RECT 14.581000  17.999000 16.330000  18.070000 ;
      RECT 14.596000  48.095000 29.845000  48.165000 ;
      RECT 14.596000  48.095000 29.845000  48.165000 ;
      RECT 14.601000  38.435000 16.069000  38.505000 ;
      RECT 14.616000  40.200000 29.845000  40.270000 ;
      RECT 14.616000  40.200000 29.845000  40.270000 ;
      RECT 14.651000   6.410000 16.815000   6.480000 ;
      RECT 14.651000   6.410000 16.815000   6.480000 ;
      RECT 14.651000  18.070000 16.330000  18.140000 ;
      RECT 14.666000  48.165000 29.845000  48.235000 ;
      RECT 14.666000  48.165000 29.845000  48.235000 ;
      RECT 14.671000  38.365000 16.139000  38.435000 ;
      RECT 14.721000   6.480000 16.815000   6.550000 ;
      RECT 14.721000   6.480000 16.815000   6.550000 ;
      RECT 14.721000  18.140000 16.330000  18.210000 ;
      RECT 14.731000   6.550000 16.815000   6.560000 ;
      RECT 14.731000   6.550000 16.815000   6.560000 ;
      RECT 14.736000  48.235000 29.845000  48.305000 ;
      RECT 14.736000  48.235000 29.845000  48.305000 ;
      RECT 14.741000  38.295000 16.209000  38.365000 ;
      RECT 14.750000  48.517000 29.985000  51.372000 ;
      RECT 14.750000  51.372000 29.567000  51.790000 ;
      RECT 14.750000  51.790000 24.535000  53.197000 ;
      RECT 14.750000  53.197000 24.535000  56.897000 ;
      RECT 14.750000  56.897000 24.212000  57.220000 ;
      RECT 14.750000  57.220000 22.940000  57.767000 ;
      RECT 14.750000  57.767000 22.940000  57.780000 ;
      RECT 14.763000  57.780000 76.775000  57.992000 ;
      RECT 14.791000  18.210000 16.330000  18.280000 ;
      RECT 14.801000   6.559000 16.744000   6.630000 ;
      RECT 14.801000   6.559000 16.744000   6.630000 ;
      RECT 14.806000  48.305000 29.845000  48.375000 ;
      RECT 14.806000  48.305000 29.845000  48.375000 ;
      RECT 14.811000  38.225000 16.279000  38.295000 ;
      RECT 14.861000  18.280000 16.330000  18.350000 ;
      RECT 14.871000   6.630000 16.674000   6.700000 ;
      RECT 14.871000   6.630000 16.674000   6.700000 ;
      RECT 14.876000  48.375000 29.845000  48.445000 ;
      RECT 14.876000  48.375000 29.845000  48.445000 ;
      RECT 14.881000  38.155000 16.349000  38.225000 ;
      RECT 14.890000  48.459000 29.845000  51.314000 ;
      RECT 14.890000  51.314000 29.774000  51.385000 ;
      RECT 14.890000  51.314000 29.774000  51.385000 ;
      RECT 14.890000  51.385000 29.704000  51.455000 ;
      RECT 14.890000  51.385000 29.704000  51.455000 ;
      RECT 14.890000  51.455000 29.634000  51.525000 ;
      RECT 14.890000  51.455000 29.634000  51.525000 ;
      RECT 14.890000  51.525000 29.564000  51.595000 ;
      RECT 14.890000  51.525000 29.564000  51.595000 ;
      RECT 14.890000  51.595000 29.509000  51.650000 ;
      RECT 14.890000  51.595000 29.509000  51.650000 ;
      RECT 14.890000  51.650000 24.395000  56.839000 ;
      RECT 14.890000  51.650000 25.814000  51.720000 ;
      RECT 14.890000  51.650000 25.814000  51.720000 ;
      RECT 14.890000  51.720000 25.744000  51.790000 ;
      RECT 14.890000  51.720000 25.744000  51.790000 ;
      RECT 14.890000  51.790000 25.674000  51.860000 ;
      RECT 14.890000  51.790000 25.674000  51.860000 ;
      RECT 14.890000  51.860000 25.604000  51.930000 ;
      RECT 14.890000  51.860000 25.604000  51.930000 ;
      RECT 14.890000  51.930000 25.534000  52.000000 ;
      RECT 14.890000  51.930000 25.534000  52.000000 ;
      RECT 14.890000  52.000000 25.464000  52.070000 ;
      RECT 14.890000  52.000000 25.464000  52.070000 ;
      RECT 14.890000  52.070000 25.394000  52.140000 ;
      RECT 14.890000  52.070000 25.394000  52.140000 ;
      RECT 14.890000  52.140000 25.324000  52.210000 ;
      RECT 14.890000  52.140000 25.324000  52.210000 ;
      RECT 14.890000  52.210000 25.254000  52.280000 ;
      RECT 14.890000  52.210000 25.254000  52.280000 ;
      RECT 14.890000  52.280000 25.184000  52.350000 ;
      RECT 14.890000  52.280000 25.184000  52.350000 ;
      RECT 14.890000  52.350000 25.114000  52.420000 ;
      RECT 14.890000  52.350000 25.114000  52.420000 ;
      RECT 14.890000  52.420000 25.044000  52.490000 ;
      RECT 14.890000  52.420000 25.044000  52.490000 ;
      RECT 14.890000  52.490000 24.974000  52.560000 ;
      RECT 14.890000  52.490000 24.974000  52.560000 ;
      RECT 14.890000  52.560000 24.904000  52.630000 ;
      RECT 14.890000  52.560000 24.904000  52.630000 ;
      RECT 14.890000  52.630000 24.834000  52.700000 ;
      RECT 14.890000  52.630000 24.834000  52.700000 ;
      RECT 14.890000  52.700000 24.764000  52.770000 ;
      RECT 14.890000  52.700000 24.764000  52.770000 ;
      RECT 14.890000  52.770000 24.694000  52.840000 ;
      RECT 14.890000  52.770000 24.694000  52.840000 ;
      RECT 14.890000  52.840000 24.624000  52.910000 ;
      RECT 14.890000  52.840000 24.624000  52.910000 ;
      RECT 14.890000  52.910000 24.554000  52.980000 ;
      RECT 14.890000  52.910000 24.554000  52.980000 ;
      RECT 14.890000  52.980000 24.484000  53.050000 ;
      RECT 14.890000  52.980000 24.484000  53.050000 ;
      RECT 14.890000  53.050000 24.414000  53.120000 ;
      RECT 14.890000  53.050000 24.414000  53.120000 ;
      RECT 14.890000  53.120000 24.394000  53.140000 ;
      RECT 14.890000  53.120000 24.394000  53.140000 ;
      RECT 14.890000  53.139000 24.395000  56.839000 ;
      RECT 14.890000  56.839000 24.324000  56.910000 ;
      RECT 14.890000  56.839000 24.324000  56.910000 ;
      RECT 14.890000  56.910000 24.254000  56.980000 ;
      RECT 14.890000  56.910000 24.254000  56.980000 ;
      RECT 14.890000  56.980000 24.184000  57.050000 ;
      RECT 14.890000  56.980000 24.184000  57.050000 ;
      RECT 14.890000  57.050000 24.154000  57.080000 ;
      RECT 14.890000  57.050000 24.154000  57.080000 ;
      RECT 14.890000  57.080000 22.800000  57.709000 ;
      RECT 14.891000  48.445000 29.845000  48.460000 ;
      RECT 14.891000  48.445000 29.845000  48.460000 ;
      RECT 14.931000  18.350000 16.330000  18.420000 ;
      RECT 14.941000   6.700000 16.604000   6.770000 ;
      RECT 14.941000   6.700000 16.604000   6.770000 ;
      RECT 14.951000  38.085000 16.419000  38.155000 ;
      RECT 14.961000  57.709000 22.800000  57.780000 ;
      RECT 14.961000  57.709000 22.800000  57.780000 ;
      RECT 14.975000  57.992000 76.775000  58.450000 ;
      RECT 15.001000  18.420000 16.330000  18.490000 ;
      RECT 15.011000   6.770000 16.534000   6.840000 ;
      RECT 15.011000   6.770000 16.534000   6.840000 ;
      RECT 15.021000  38.015000 16.489000  38.085000 ;
      RECT 15.031000  57.780000 22.800000  57.850000 ;
      RECT 15.031000  57.780000 22.800000  57.850000 ;
      RECT 15.071000  18.490000 16.330000  18.560000 ;
      RECT 15.081000   6.840000 16.464000   6.910000 ;
      RECT 15.081000   6.840000 16.464000   6.910000 ;
      RECT 15.091000  37.945000 16.559000  38.015000 ;
      RECT 15.101000  57.850000 22.800000  57.920000 ;
      RECT 15.101000  57.850000 22.800000  57.920000 ;
      RECT 15.106000  57.920000 76.635000  57.925000 ;
      RECT 15.106000  57.920000 76.635000  57.925000 ;
      RECT 15.111000  57.925000 76.635000  57.930000 ;
      RECT 15.111000  57.925000 76.635000  57.930000 ;
      RECT 15.115000  57.920000 76.635000  73.499000 ;
      RECT 15.115000  57.920000 76.635000  73.499000 ;
      RECT 15.115000  57.920000 76.635000  73.499000 ;
      RECT 15.115000  57.920000 76.635000  73.499000 ;
      RECT 15.115000  57.934000 76.635000  58.590000 ;
      RECT 15.116000  57.930000 76.635000  57.935000 ;
      RECT 15.116000  57.930000 76.635000  57.935000 ;
      RECT 15.141000  18.560000 16.330000  18.630000 ;
      RECT 15.151000   6.910000 16.394000   6.980000 ;
      RECT 15.151000   6.910000 16.394000   6.980000 ;
      RECT 15.161000  37.875000 16.629000  37.945000 ;
      RECT 15.211000  18.630000 16.330000  18.700000 ;
      RECT 15.216000   6.980000 16.329000   7.045000 ;
      RECT 15.216000   6.980000 16.329000   7.045000 ;
      RECT 15.231000  37.805000 16.699000  37.875000 ;
      RECT 15.281000  18.700000 16.330000  18.770000 ;
      RECT 15.301000  37.735000 16.769000  37.805000 ;
      RECT 15.351000  18.770000 16.330000  18.840000 ;
      RECT 15.370000  32.128000 16.225000  34.378000 ;
      RECT 15.370000  34.378000 17.435000  35.588000 ;
      RECT 15.370000  35.588000 17.435000  37.337000 ;
      RECT 15.370000  37.337000 17.304000  37.468000 ;
      RECT 15.371000  37.665000 16.839000  37.735000 ;
      RECT 15.421000  18.840000 16.330000  18.910000 ;
      RECT 15.441000  37.595000 16.909000  37.665000 ;
      RECT 15.491000  18.910000 16.330000  18.980000 ;
      RECT 15.510000  32.186000 16.085000  34.436000 ;
      RECT 15.510000  34.436000 16.085000  34.505000 ;
      RECT 15.510000  34.505000 16.154000  34.575000 ;
      RECT 15.510000  34.575000 16.224000  34.645000 ;
      RECT 15.510000  34.645000 16.294000  34.715000 ;
      RECT 15.510000  34.715000 16.364000  34.785000 ;
      RECT 15.510000  34.785000 16.434000  34.855000 ;
      RECT 15.510000  34.855000 16.504000  34.925000 ;
      RECT 15.510000  34.925000 16.574000  34.995000 ;
      RECT 15.510000  34.995000 16.644000  35.065000 ;
      RECT 15.510000  35.065000 16.714000  35.135000 ;
      RECT 15.510000  35.135000 16.784000  35.205000 ;
      RECT 15.510000  35.205000 16.854000  35.275000 ;
      RECT 15.510000  35.275000 16.924000  35.345000 ;
      RECT 15.510000  35.345000 16.994000  35.415000 ;
      RECT 15.510000  35.415000 17.064000  35.485000 ;
      RECT 15.510000  35.485000 17.134000  35.555000 ;
      RECT 15.510000  35.555000 17.204000  35.625000 ;
      RECT 15.510000  35.625000 17.274000  35.645000 ;
      RECT 15.510000  35.646000 17.295000  37.279000 ;
      RECT 15.510000  37.279000 17.224000  37.350000 ;
      RECT 15.510000  37.350000 17.154000  37.420000 ;
      RECT 15.510000  37.420000 17.084000  37.490000 ;
      RECT 15.510000  37.490000 17.049000  37.525000 ;
      RECT 15.510000  37.526000 16.979000  37.595000 ;
      RECT 15.561000  18.980000 16.330000  19.050000 ;
      RECT 15.576000  32.120000 16.085000  32.185000 ;
      RECT 15.591000  40.145000 29.845000  40.200000 ;
      RECT 15.591000  40.145000 29.845000  40.200000 ;
      RECT 15.631000  19.050000 16.330000  19.120000 ;
      RECT 15.646000  32.050000 16.085000  32.120000 ;
      RECT 15.661000  40.075000 29.845000  40.145000 ;
      RECT 15.661000  40.075000 29.845000  40.145000 ;
      RECT 15.701000  19.120000 16.330000  19.190000 ;
      RECT 15.716000  31.980000 16.085000  32.050000 ;
      RECT 15.731000  40.005000 29.845000  40.075000 ;
      RECT 15.731000  40.005000 29.845000  40.075000 ;
      RECT 15.771000  19.190000 16.330000  19.260000 ;
      RECT 15.785000  19.472000 16.470000  31.257000 ;
      RECT 15.785000  31.257000 16.225000  31.502000 ;
      RECT 15.785000  31.502000 16.225000  31.713000 ;
      RECT 15.785000  31.713000 16.225000  32.128000 ;
      RECT 15.786000  31.910000 16.085000  31.980000 ;
      RECT 15.801000  39.935000 29.845000  40.005000 ;
      RECT 15.801000  39.935000 29.845000  40.005000 ;
      RECT 15.841000  19.260000 16.330000  19.330000 ;
      RECT 15.856000  31.840000 16.085000  31.910000 ;
      RECT 15.871000  39.865000 29.845000  39.935000 ;
      RECT 15.871000  39.865000 29.845000  39.935000 ;
      RECT 15.911000  19.330000 16.330000  19.400000 ;
      RECT 15.925000  19.414000 16.330000  31.199000 ;
      RECT 15.925000  31.199000 16.259000  31.270000 ;
      RECT 15.925000  31.270000 16.189000  31.340000 ;
      RECT 15.925000  31.340000 16.119000  31.410000 ;
      RECT 15.925000  31.410000 16.084000  31.445000 ;
      RECT 15.925000  31.444000 16.085000  31.771000 ;
      RECT 15.925000  31.771000 16.085000  31.840000 ;
      RECT 15.926000  19.400000 16.330000  19.415000 ;
      RECT 15.941000  39.795000 29.845000  39.865000 ;
      RECT 15.941000  39.795000 29.845000  39.865000 ;
      RECT 16.011000  39.725000 29.845000  39.795000 ;
      RECT 16.011000  39.725000 29.845000  39.795000 ;
      RECT 16.081000  39.655000 29.845000  39.725000 ;
      RECT 16.081000  39.655000 29.845000  39.725000 ;
      RECT 16.151000  39.585000 29.845000  39.655000 ;
      RECT 16.151000  39.585000 29.845000  39.655000 ;
      RECT 16.221000  39.515000 29.845000  39.585000 ;
      RECT 16.221000  39.515000 29.845000  39.585000 ;
      RECT 16.291000  39.445000 29.845000  39.515000 ;
      RECT 16.291000  39.445000 29.845000  39.515000 ;
      RECT 16.361000  39.375000 29.845000  39.445000 ;
      RECT 16.361000  39.375000 29.845000  39.445000 ;
      RECT 16.431000  39.305000 29.845000  39.375000 ;
      RECT 16.431000  39.305000 29.845000  39.375000 ;
      RECT 16.443000  39.095000 29.985000  40.060000 ;
      RECT 16.501000  39.235000 29.845000  39.305000 ;
      RECT 16.501000  39.235000 29.845000  39.305000 ;
      RECT 16.551000  39.185000 22.815000  39.235000 ;
      RECT 16.551000  39.185000 22.815000  39.235000 ;
      RECT 16.621000  39.115000 22.815000  39.185000 ;
      RECT 16.621000  39.115000 22.815000  39.185000 ;
      RECT 16.691000  39.045000 22.815000  39.115000 ;
      RECT 16.691000  39.045000 22.815000  39.115000 ;
      RECT 16.710000   0.000000 22.215000   2.152000 ;
      RECT 16.710000   2.152000 22.215000   2.937000 ;
      RECT 16.761000  38.975000 22.815000  39.045000 ;
      RECT 16.761000  38.975000 22.815000  39.045000 ;
      RECT 16.765000  31.728000 23.335000  34.152000 ;
      RECT 16.765000  34.152000 23.335000  35.362000 ;
      RECT 16.831000  38.905000 22.815000  38.975000 ;
      RECT 16.831000  38.905000 22.815000  38.975000 ;
      RECT 16.850000   0.000000 22.075000   2.094000 ;
      RECT 16.901000  38.835000 22.815000  38.905000 ;
      RECT 16.901000  38.835000 22.815000  38.905000 ;
      RECT 16.905000  31.786000 23.195000  34.094000 ;
      RECT 16.921000   2.094000 22.075000   2.165000 ;
      RECT 16.921000   2.094000 22.075000   2.165000 ;
      RECT 16.941000  31.750000 23.195000  31.785000 ;
      RECT 16.941000  31.750000 23.195000  31.785000 ;
      RECT 16.971000  38.765000 22.815000  38.835000 ;
      RECT 16.971000  38.765000 22.815000  38.835000 ;
      RECT 16.976000  34.094000 23.195000  34.165000 ;
      RECT 16.976000  34.094000 23.195000  34.165000 ;
      RECT 16.983000  38.555000 22.955000  39.095000 ;
      RECT 16.991000   2.165000 22.075000   2.235000 ;
      RECT 16.991000   2.165000 22.075000   2.235000 ;
      RECT 17.010000   7.328000 22.625000  14.543000 ;
      RECT 17.010000  14.543000 23.515000  15.433000 ;
      RECT 17.010000  15.433000 23.515000  24.942000 ;
      RECT 17.010000  24.942000 23.335000  25.122000 ;
      RECT 17.010000  25.122000 23.335000  31.483000 ;
      RECT 17.010000  31.483000 23.335000  31.728000 ;
      RECT 17.011000  31.680000 23.195000  31.750000 ;
      RECT 17.011000  31.680000 23.195000  31.750000 ;
      RECT 17.041000  38.695000 22.815000  38.765000 ;
      RECT 17.041000  38.695000 22.815000  38.765000 ;
      RECT 17.046000  34.165000 23.195000  34.235000 ;
      RECT 17.046000  34.165000 23.195000  34.235000 ;
      RECT 17.061000   2.235000 22.075000   2.305000 ;
      RECT 17.061000   2.235000 22.075000   2.305000 ;
      RECT 17.081000  31.610000 23.195000  31.680000 ;
      RECT 17.081000  31.610000 23.195000  31.680000 ;
      RECT 17.111000  38.625000 22.815000  38.695000 ;
      RECT 17.111000  38.625000 22.815000  38.695000 ;
      RECT 17.116000  34.235000 23.195000  34.305000 ;
      RECT 17.116000  34.235000 23.195000  34.305000 ;
      RECT 17.131000   2.305000 22.075000   2.375000 ;
      RECT 17.131000   2.305000 22.075000   2.375000 ;
      RECT 17.150000   7.386000 22.485000  14.601000 ;
      RECT 17.150000   7.386000 22.485000  15.491000 ;
      RECT 17.150000  14.601000 22.485000  14.670000 ;
      RECT 17.150000  14.601000 22.485000  14.670000 ;
      RECT 17.150000  14.670000 22.554000  14.740000 ;
      RECT 17.150000  14.670000 22.554000  14.740000 ;
      RECT 17.150000  14.740000 22.624000  14.810000 ;
      RECT 17.150000  14.740000 22.624000  14.810000 ;
      RECT 17.150000  14.810000 22.694000  14.880000 ;
      RECT 17.150000  14.810000 22.694000  14.880000 ;
      RECT 17.150000  14.880000 22.764000  14.950000 ;
      RECT 17.150000  14.880000 22.764000  14.950000 ;
      RECT 17.150000  14.950000 22.834000  15.020000 ;
      RECT 17.150000  14.950000 22.834000  15.020000 ;
      RECT 17.150000  15.020000 22.904000  15.090000 ;
      RECT 17.150000  15.020000 22.904000  15.090000 ;
      RECT 17.150000  15.090000 22.974000  15.160000 ;
      RECT 17.150000  15.090000 22.974000  15.160000 ;
      RECT 17.150000  15.160000 23.044000  15.230000 ;
      RECT 17.150000  15.160000 23.044000  15.230000 ;
      RECT 17.150000  15.230000 23.114000  15.300000 ;
      RECT 17.150000  15.230000 23.114000  15.300000 ;
      RECT 17.150000  15.300000 23.184000  15.370000 ;
      RECT 17.150000  15.300000 23.184000  15.370000 ;
      RECT 17.150000  15.370000 23.254000  15.440000 ;
      RECT 17.150000  15.370000 23.254000  15.440000 ;
      RECT 17.150000  15.440000 23.324000  15.490000 ;
      RECT 17.150000  15.440000 23.324000  15.490000 ;
      RECT 17.150000  15.491000 23.375000  24.884000 ;
      RECT 17.150000  24.884000 23.304000  24.955000 ;
      RECT 17.150000  24.884000 23.304000  24.955000 ;
      RECT 17.150000  24.955000 23.234000  25.025000 ;
      RECT 17.150000  24.955000 23.234000  25.025000 ;
      RECT 17.150000  25.025000 23.194000  25.065000 ;
      RECT 17.150000  25.025000 23.194000  25.065000 ;
      RECT 17.150000  25.064000 23.195000  31.541000 ;
      RECT 17.150000  31.541000 23.195000  31.610000 ;
      RECT 17.150000  31.541000 23.195000  31.610000 ;
      RECT 17.166000   7.370000 22.485000   7.385000 ;
      RECT 17.166000   7.370000 22.485000   7.385000 ;
      RECT 17.181000  38.357000 23.137000  38.555000 ;
      RECT 17.181000  38.555000 22.815000  38.625000 ;
      RECT 17.181000  38.555000 22.815000  38.625000 ;
      RECT 17.186000  34.305000 23.195000  34.375000 ;
      RECT 17.186000  34.305000 23.195000  34.375000 ;
      RECT 17.201000   2.375000 22.075000   2.445000 ;
      RECT 17.201000   2.375000 22.075000   2.445000 ;
      RECT 17.236000   7.300000 22.485000   7.370000 ;
      RECT 17.236000   7.300000 22.485000   7.370000 ;
      RECT 17.251000  38.485000 22.815000  38.555000 ;
      RECT 17.251000  38.485000 22.815000  38.555000 ;
      RECT 17.256000  34.375000 23.195000  34.445000 ;
      RECT 17.256000  34.375000 23.195000  34.445000 ;
      RECT 17.271000   2.445000 22.075000   2.515000 ;
      RECT 17.271000   2.445000 22.075000   2.515000 ;
      RECT 17.306000   7.230000 22.485000   7.300000 ;
      RECT 17.306000   7.230000 22.485000   7.300000 ;
      RECT 17.321000  38.415000 22.815000  38.485000 ;
      RECT 17.321000  38.415000 22.815000  38.485000 ;
      RECT 17.326000  34.445000 23.195000  34.515000 ;
      RECT 17.326000  34.445000 23.195000  34.515000 ;
      RECT 17.341000   2.515000 22.075000   2.585000 ;
      RECT 17.341000   2.515000 22.075000   2.585000 ;
      RECT 17.376000   7.160000 22.485000   7.230000 ;
      RECT 17.376000   7.160000 22.485000   7.230000 ;
      RECT 17.381000  38.355000 23.079000  38.415000 ;
      RECT 17.381000  38.355000 23.079000  38.415000 ;
      RECT 17.396000  34.515000 23.195000  34.585000 ;
      RECT 17.396000  34.515000 23.195000  34.585000 ;
      RECT 17.411000   2.585000 22.075000   2.655000 ;
      RECT 17.411000   2.585000 22.075000   2.655000 ;
      RECT 17.437000  38.299000 23.139000  38.355000 ;
      RECT 17.437000  38.299000 23.139000  38.355000 ;
      RECT 17.445000   6.893000 22.625000   7.328000 ;
      RECT 17.446000   7.090000 22.485000   7.160000 ;
      RECT 17.446000   7.090000 22.485000   7.160000 ;
      RECT 17.466000  34.585000 23.195000  34.655000 ;
      RECT 17.466000  34.585000 23.195000  34.655000 ;
      RECT 17.481000   2.655000 22.075000   2.725000 ;
      RECT 17.481000   2.655000 22.075000   2.725000 ;
      RECT 17.486000  38.250000 23.195000  38.300000 ;
      RECT 17.486000  38.250000 23.195000  38.300000 ;
      RECT 17.495000   2.937000 22.215000   6.483000 ;
      RECT 17.495000   6.483000 22.575000   6.843000 ;
      RECT 17.495000   6.843000 22.625000   6.893000 ;
      RECT 17.516000   7.020000 22.485000   7.090000 ;
      RECT 17.516000   7.020000 22.485000   7.090000 ;
      RECT 17.536000  34.655000 23.195000  34.725000 ;
      RECT 17.536000  34.655000 23.195000  34.725000 ;
      RECT 17.551000   2.725000 22.075000   2.795000 ;
      RECT 17.551000   2.725000 22.075000   2.795000 ;
      RECT 17.556000  38.180000 23.195000  38.250000 ;
      RECT 17.556000  38.180000 23.195000  38.250000 ;
      RECT 17.585000   6.951000 22.485000   7.020000 ;
      RECT 17.585000   6.951000 22.485000   7.020000 ;
      RECT 17.606000  34.725000 23.195000  34.795000 ;
      RECT 17.606000  34.725000 23.195000  34.795000 ;
      RECT 17.611000   6.925000 22.459000   6.950000 ;
      RECT 17.611000   6.925000 22.459000   6.950000 ;
      RECT 17.621000   2.795000 22.075000   2.865000 ;
      RECT 17.621000   2.795000 22.075000   2.865000 ;
      RECT 17.626000  38.110000 23.195000  38.180000 ;
      RECT 17.626000  38.110000 23.195000  38.180000 ;
      RECT 17.635000   0.000000 22.075000   6.541000 ;
      RECT 17.635000   0.000000 22.075000   6.541000 ;
      RECT 17.635000   2.879000 22.075000   6.541000 ;
      RECT 17.635000   2.879000 22.075000   6.901000 ;
      RECT 17.635000   2.879000 22.075000   6.901000 ;
      RECT 17.635000   2.879000 22.075000   6.901000 ;
      RECT 17.635000   2.879000 22.075000   6.901000 ;
      RECT 17.635000   6.541000 22.075000   6.610000 ;
      RECT 17.635000   6.541000 22.075000   6.610000 ;
      RECT 17.635000   6.610000 22.144000   6.680000 ;
      RECT 17.635000   6.610000 22.144000   6.680000 ;
      RECT 17.635000   6.680000 22.214000   6.750000 ;
      RECT 17.635000   6.680000 22.214000   6.750000 ;
      RECT 17.635000   6.750000 22.284000   6.820000 ;
      RECT 17.635000   6.750000 22.284000   6.820000 ;
      RECT 17.635000   6.820000 22.354000   6.890000 ;
      RECT 17.635000   6.820000 22.354000   6.890000 ;
      RECT 17.635000   6.890000 22.424000   6.900000 ;
      RECT 17.635000   6.890000 22.424000   6.900000 ;
      RECT 17.635000   6.901000 22.435000   6.925000 ;
      RECT 17.635000   6.901000 22.435000   6.925000 ;
      RECT 17.636000   2.865000 22.075000   2.880000 ;
      RECT 17.636000   2.865000 22.075000   2.880000 ;
      RECT 17.676000  34.795000 23.195000  34.865000 ;
      RECT 17.676000  34.795000 23.195000  34.865000 ;
      RECT 17.696000  38.040000 23.195000  38.110000 ;
      RECT 17.696000  38.040000 23.195000  38.110000 ;
      RECT 17.746000  34.865000 23.195000  34.935000 ;
      RECT 17.746000  34.865000 23.195000  34.935000 ;
      RECT 17.766000  37.970000 23.195000  38.040000 ;
      RECT 17.766000  37.970000 23.195000  38.040000 ;
      RECT 17.816000  34.935000 23.195000  35.005000 ;
      RECT 17.816000  34.935000 23.195000  35.005000 ;
      RECT 17.836000  37.900000 23.195000  37.970000 ;
      RECT 17.836000  37.900000 23.195000  37.970000 ;
      RECT 17.886000  35.005000 23.195000  35.075000 ;
      RECT 17.886000  35.005000 23.195000  35.075000 ;
      RECT 17.906000  37.830000 23.195000  37.900000 ;
      RECT 17.906000  37.830000 23.195000  37.900000 ;
      RECT 17.956000  35.075000 23.195000  35.145000 ;
      RECT 17.956000  35.075000 23.195000  35.145000 ;
      RECT 17.975000  35.362000 23.335000  37.563000 ;
      RECT 17.975000  37.563000 23.335000  38.357000 ;
      RECT 17.976000  37.760000 23.195000  37.830000 ;
      RECT 17.976000  37.760000 23.195000  37.830000 ;
      RECT 18.026000  35.145000 23.195000  35.215000 ;
      RECT 18.026000  35.145000 23.195000  35.215000 ;
      RECT 18.046000  37.690000 23.195000  37.760000 ;
      RECT 18.046000  37.690000 23.195000  37.760000 ;
      RECT 18.096000  35.215000 23.195000  35.285000 ;
      RECT 18.096000  35.215000 23.195000  35.285000 ;
      RECT 18.115000  31.541000 23.195000  37.621000 ;
      RECT 18.115000  35.304000 23.195000  37.621000 ;
      RECT 18.115000  37.621000 23.195000  37.690000 ;
      RECT 18.115000  37.621000 23.195000  37.690000 ;
      RECT 18.116000  35.285000 23.195000  35.305000 ;
      RECT 18.116000  35.285000 23.195000  35.305000 ;
      RECT 22.755000   0.000000 26.460000   1.835000 ;
      RECT 22.755000   1.835000 28.350000   4.128000 ;
      RECT 22.755000   4.128000 29.070000   4.848000 ;
      RECT 22.755000   4.848000 29.070000   6.257000 ;
      RECT 22.755000   6.257000 29.070000   6.667000 ;
      RECT 22.895000   0.000000 26.320000   1.975000 ;
      RECT 22.895000   0.000000 26.320000   4.186000 ;
      RECT 22.895000   0.000000 26.320000   6.199000 ;
      RECT 22.895000   0.000000 26.320000   6.199000 ;
      RECT 22.895000   0.000000 26.320000   6.199000 ;
      RECT 22.895000   1.975000 28.210000   4.186000 ;
      RECT 22.895000   1.975000 28.210000   6.199000 ;
      RECT 22.895000   1.975000 28.210000   6.199000 ;
      RECT 22.895000   1.975000 28.210000   6.199000 ;
      RECT 22.895000   1.975000 28.210000   6.199000 ;
      RECT 22.895000   1.975000 28.210000   6.199000 ;
      RECT 22.895000   4.186000 28.210000   4.255000 ;
      RECT 22.895000   4.186000 28.210000   4.255000 ;
      RECT 22.895000   4.255000 28.279000   4.325000 ;
      RECT 22.895000   4.255000 28.279000   4.325000 ;
      RECT 22.895000   4.325000 28.349000   4.395000 ;
      RECT 22.895000   4.325000 28.349000   4.395000 ;
      RECT 22.895000   4.395000 28.419000   4.465000 ;
      RECT 22.895000   4.395000 28.419000   4.465000 ;
      RECT 22.895000   4.465000 28.489000   4.535000 ;
      RECT 22.895000   4.465000 28.489000   4.535000 ;
      RECT 22.895000   4.535000 28.559000   4.605000 ;
      RECT 22.895000   4.535000 28.559000   4.605000 ;
      RECT 22.895000   4.605000 28.629000   4.675000 ;
      RECT 22.895000   4.605000 28.629000   4.675000 ;
      RECT 22.895000   4.675000 28.699000   4.745000 ;
      RECT 22.895000   4.675000 28.699000   4.745000 ;
      RECT 22.895000   4.745000 28.769000   4.815000 ;
      RECT 22.895000   4.745000 28.769000   4.815000 ;
      RECT 22.895000   4.815000 28.839000   4.885000 ;
      RECT 22.895000   4.815000 28.839000   4.885000 ;
      RECT 22.895000   4.885000 28.909000   4.905000 ;
      RECT 22.895000   4.885000 28.909000   4.905000 ;
      RECT 22.895000   4.906000 28.930000   6.199000 ;
      RECT 22.966000   6.199000 28.930000   6.270000 ;
      RECT 22.966000   6.199000 28.930000   6.270000 ;
      RECT 23.036000   6.270000 28.930000   6.340000 ;
      RECT 23.036000   6.270000 28.930000   6.340000 ;
      RECT 23.106000   6.340000 28.930000   6.410000 ;
      RECT 23.106000   6.340000 28.930000   6.410000 ;
      RECT 23.165000   6.667000 29.070000   6.920000 ;
      RECT 23.165000   6.920000 31.550000  14.317000 ;
      RECT 23.165000  14.317000 31.550000  15.207000 ;
      RECT 23.176000   6.410000 28.930000   6.480000 ;
      RECT 23.176000   6.410000 28.930000   6.480000 ;
      RECT 23.246000   6.480000 28.930000   6.550000 ;
      RECT 23.246000   6.480000 28.930000   6.550000 ;
      RECT 23.305000   6.609000 28.930000   7.060000 ;
      RECT 23.305000   7.060000 31.410000  14.259000 ;
      RECT 23.306000   6.550000 28.930000   6.610000 ;
      RECT 23.306000   6.550000 28.930000   6.610000 ;
      RECT 23.376000  14.259000 31.410000  14.330000 ;
      RECT 23.376000  14.259000 31.410000  14.330000 ;
      RECT 23.446000  14.330000 31.410000  14.400000 ;
      RECT 23.446000  14.330000 31.410000  14.400000 ;
      RECT 23.516000  14.400000 31.410000  14.470000 ;
      RECT 23.516000  14.400000 31.410000  14.470000 ;
      RECT 23.586000  14.470000 31.410000  14.540000 ;
      RECT 23.586000  14.470000 31.410000  14.540000 ;
      RECT 23.656000  14.540000 31.410000  14.610000 ;
      RECT 23.656000  14.540000 31.410000  14.610000 ;
      RECT 23.726000  14.610000 31.410000  14.680000 ;
      RECT 23.726000  14.610000 31.410000  14.680000 ;
      RECT 23.796000  14.680000 31.410000  14.750000 ;
      RECT 23.796000  14.680000 31.410000  14.750000 ;
      RECT 23.866000  14.750000 31.410000  14.820000 ;
      RECT 23.866000  14.750000 31.410000  14.820000 ;
      RECT 23.875000  25.348000 29.985000  36.513000 ;
      RECT 23.875000  36.513000 30.250000  36.778000 ;
      RECT 23.875000  36.778000 30.250000  37.687000 ;
      RECT 23.875000  37.687000 29.985000  37.952000 ;
      RECT 23.875000  37.952000 29.985000  39.095000 ;
      RECT 23.936000  14.820000 31.410000  14.890000 ;
      RECT 23.936000  14.820000 31.410000  14.890000 ;
      RECT 24.006000  14.890000 31.410000  14.960000 ;
      RECT 24.006000  14.890000 31.410000  14.960000 ;
      RECT 24.015000  25.406000 29.845000  37.629000 ;
      RECT 24.015000  36.571000 29.845000  36.640000 ;
      RECT 24.015000  36.571000 29.845000  36.640000 ;
      RECT 24.015000  36.640000 29.914000  36.710000 ;
      RECT 24.015000  36.640000 29.914000  36.710000 ;
      RECT 24.015000  36.710000 29.984000  36.780000 ;
      RECT 24.015000  36.710000 29.984000  36.780000 ;
      RECT 24.015000  36.780000 30.054000  36.835000 ;
      RECT 24.015000  36.780000 30.054000  36.835000 ;
      RECT 24.015000  36.836000 30.110000  37.246000 ;
      RECT 24.015000  37.246000 30.110000  37.629000 ;
      RECT 24.015000  37.629000 30.039000  37.700000 ;
      RECT 24.015000  37.629000 30.039000  37.700000 ;
      RECT 24.015000  37.700000 29.969000  37.770000 ;
      RECT 24.015000  37.700000 29.969000  37.770000 ;
      RECT 24.015000  37.770000 29.899000  37.840000 ;
      RECT 24.015000  37.770000 29.899000  37.840000 ;
      RECT 24.015000  37.840000 29.844000  37.895000 ;
      RECT 24.015000  37.840000 29.844000  37.895000 ;
      RECT 24.015000  37.894000 29.845000  39.235000 ;
      RECT 24.055000  15.207000 31.550000  16.007000 ;
      RECT 24.055000  16.007000 29.985000  17.572000 ;
      RECT 24.055000  17.572000 29.985000  25.168000 ;
      RECT 24.055000  25.168000 29.985000  25.348000 ;
      RECT 24.056000  25.365000 29.845000  25.405000 ;
      RECT 24.056000  25.365000 29.845000  25.405000 ;
      RECT 24.076000  14.960000 31.410000  15.030000 ;
      RECT 24.076000  14.960000 31.410000  15.030000 ;
      RECT 24.126000  25.295000 29.845000  25.365000 ;
      RECT 24.126000  25.295000 29.845000  25.365000 ;
      RECT 24.146000  15.030000 31.410000  15.100000 ;
      RECT 24.146000  15.030000 31.410000  15.100000 ;
      RECT 24.195000  15.149000 31.410000  15.949000 ;
      RECT 24.195000  15.949000 29.845000  25.226000 ;
      RECT 24.195000  15.949000 31.339000  16.020000 ;
      RECT 24.195000  15.949000 31.339000  16.020000 ;
      RECT 24.195000  16.020000 31.269000  16.090000 ;
      RECT 24.195000  16.020000 31.269000  16.090000 ;
      RECT 24.195000  16.090000 31.199000  16.160000 ;
      RECT 24.195000  16.090000 31.199000  16.160000 ;
      RECT 24.195000  16.160000 31.129000  16.230000 ;
      RECT 24.195000  16.160000 31.129000  16.230000 ;
      RECT 24.195000  16.230000 31.059000  16.300000 ;
      RECT 24.195000  16.230000 31.059000  16.300000 ;
      RECT 24.195000  16.300000 30.989000  16.370000 ;
      RECT 24.195000  16.300000 30.989000  16.370000 ;
      RECT 24.195000  16.370000 30.919000  16.440000 ;
      RECT 24.195000  16.370000 30.919000  16.440000 ;
      RECT 24.195000  16.440000 30.849000  16.510000 ;
      RECT 24.195000  16.440000 30.849000  16.510000 ;
      RECT 24.195000  16.510000 30.779000  16.580000 ;
      RECT 24.195000  16.510000 30.779000  16.580000 ;
      RECT 24.195000  16.580000 30.709000  16.650000 ;
      RECT 24.195000  16.580000 30.709000  16.650000 ;
      RECT 24.195000  16.650000 30.639000  16.720000 ;
      RECT 24.195000  16.650000 30.639000  16.720000 ;
      RECT 24.195000  16.720000 30.569000  16.790000 ;
      RECT 24.195000  16.720000 30.569000  16.790000 ;
      RECT 24.195000  16.790000 30.499000  16.860000 ;
      RECT 24.195000  16.790000 30.499000  16.860000 ;
      RECT 24.195000  16.860000 30.429000  16.930000 ;
      RECT 24.195000  16.860000 30.429000  16.930000 ;
      RECT 24.195000  16.930000 30.359000  17.000000 ;
      RECT 24.195000  16.930000 30.359000  17.000000 ;
      RECT 24.195000  17.000000 30.289000  17.070000 ;
      RECT 24.195000  17.000000 30.289000  17.070000 ;
      RECT 24.195000  17.070000 30.219000  17.140000 ;
      RECT 24.195000  17.070000 30.219000  17.140000 ;
      RECT 24.195000  17.140000 30.149000  17.210000 ;
      RECT 24.195000  17.140000 30.149000  17.210000 ;
      RECT 24.195000  17.210000 30.079000  17.280000 ;
      RECT 24.195000  17.210000 30.079000  17.280000 ;
      RECT 24.195000  17.280000 30.009000  17.350000 ;
      RECT 24.195000  17.280000 30.009000  17.350000 ;
      RECT 24.195000  17.350000 29.939000  17.420000 ;
      RECT 24.195000  17.350000 29.939000  17.420000 ;
      RECT 24.195000  17.420000 29.869000  17.490000 ;
      RECT 24.195000  17.420000 29.869000  17.490000 ;
      RECT 24.195000  17.490000 29.844000  17.515000 ;
      RECT 24.195000  17.490000 29.844000  17.515000 ;
      RECT 24.195000  17.514000 29.845000  25.226000 ;
      RECT 24.195000  25.226000 29.845000  25.295000 ;
      RECT 24.195000  25.226000 29.845000  25.295000 ;
      RECT 24.196000  15.100000 31.410000  15.150000 ;
      RECT 24.196000  15.100000 31.410000  15.150000 ;
      RECT 24.536000  57.880000 76.635000  57.920000 ;
      RECT 24.536000  57.880000 76.635000  57.920000 ;
      RECT 24.606000  57.810000 76.635000  57.880000 ;
      RECT 24.606000  57.810000 76.635000  57.880000 ;
      RECT 24.676000  57.740000 76.635000  57.810000 ;
      RECT 24.676000  57.740000 76.635000  57.810000 ;
      RECT 24.746000  57.670000 76.635000  57.740000 ;
      RECT 24.746000  57.670000 76.635000  57.740000 ;
      RECT 24.816000  57.600000 76.635000  57.670000 ;
      RECT 24.816000  57.600000 76.635000  57.670000 ;
      RECT 24.886000  57.530000 76.635000  57.600000 ;
      RECT 24.886000  57.530000 76.635000  57.600000 ;
      RECT 24.956000  57.460000 76.635000  57.530000 ;
      RECT 24.956000  57.460000 76.635000  57.530000 ;
      RECT 25.026000  57.390000 76.635000  57.460000 ;
      RECT 25.026000  57.390000 76.635000  57.460000 ;
      RECT 25.095000  53.423000 76.775000  57.123000 ;
      RECT 25.095000  57.123000 76.775000  57.780000 ;
      RECT 25.096000  57.320000 76.635000  57.390000 ;
      RECT 25.096000  57.320000 76.635000  57.390000 ;
      RECT 25.166000  57.250000 76.635000  57.320000 ;
      RECT 25.166000  57.250000 76.635000  57.320000 ;
      RECT 25.235000  53.481000 76.635000  57.181000 ;
      RECT 25.235000  53.481000 76.635000  57.920000 ;
      RECT 25.235000  53.481000 76.635000  73.499000 ;
      RECT 25.235000  57.181000 76.635000  57.250000 ;
      RECT 25.235000  57.181000 76.635000  57.250000 ;
      RECT 25.260000  53.258000 76.775000  53.423000 ;
      RECT 25.261000  53.455000 76.635000  53.480000 ;
      RECT 25.261000  53.455000 76.635000  53.480000 ;
      RECT 25.331000  53.385000 76.635000  53.455000 ;
      RECT 25.331000  53.385000 76.635000  53.455000 ;
      RECT 25.400000  53.316000 76.635000  53.385000 ;
      RECT 25.400000  53.316000 76.635000  53.385000 ;
      RECT 25.456000  53.260000 76.579000  53.315000 ;
      RECT 25.456000  53.260000 76.579000  53.315000 ;
      RECT 25.526000  53.190000 76.509000  53.260000 ;
      RECT 25.526000  53.190000 76.509000  53.260000 ;
      RECT 25.596000  53.120000 76.439000  53.190000 ;
      RECT 25.596000  53.120000 76.439000  53.190000 ;
      RECT 25.666000  53.050000 76.369000  53.120000 ;
      RECT 25.666000  53.050000 76.369000  53.120000 ;
      RECT 25.736000  52.980000 76.299000  53.050000 ;
      RECT 25.736000  52.980000 76.299000  53.050000 ;
      RECT 25.806000  52.910000 76.229000  52.980000 ;
      RECT 25.806000  52.910000 76.229000  52.980000 ;
      RECT 25.876000  52.840000 76.159000  52.910000 ;
      RECT 25.876000  52.840000 76.159000  52.910000 ;
      RECT 25.945000  52.573000 76.775000  53.258000 ;
      RECT 25.946000  52.770000 76.089000  52.840000 ;
      RECT 25.946000  52.770000 76.089000  52.840000 ;
      RECT 26.016000  52.700000 76.019000  52.770000 ;
      RECT 26.016000  52.700000 76.019000  52.770000 ;
      RECT 26.085000  52.631000 75.950000  52.700000 ;
      RECT 26.085000  52.631000 75.950000  52.700000 ;
      RECT 26.156000  52.560000 75.950000  52.630000 ;
      RECT 26.156000  52.560000 75.950000  52.630000 ;
      RECT 26.168000  52.350000 76.090000  52.573000 ;
      RECT 26.226000  52.490000 75.950000  52.560000 ;
      RECT 26.226000  52.490000 75.950000  52.560000 ;
      RECT 27.000000   0.000000 28.350000   1.835000 ;
      RECT 27.140000   0.000000 28.210000   1.975000 ;
      RECT 28.890000   0.000000 30.610000   2.323000 ;
      RECT 28.890000   2.323000 31.165000   2.878000 ;
      RECT 28.890000   2.878000 31.165000   3.902000 ;
      RECT 28.890000   3.902000 31.165000   4.503000 ;
      RECT 29.030000   0.000000 30.470000   2.381000 ;
      RECT 29.030000   2.381000 30.470000   2.450000 ;
      RECT 29.030000   2.450000 30.539000   2.520000 ;
      RECT 29.030000   2.520000 30.609000   2.590000 ;
      RECT 29.030000   2.590000 30.679000   2.660000 ;
      RECT 29.030000   2.660000 30.749000   2.730000 ;
      RECT 29.030000   2.730000 30.819000   2.800000 ;
      RECT 29.030000   2.800000 30.889000   2.870000 ;
      RECT 29.030000   2.870000 30.959000   2.935000 ;
      RECT 29.030000   2.936000 31.025000   3.844000 ;
      RECT 29.101000   3.844000 31.025000   3.915000 ;
      RECT 29.171000   3.915000 31.025000   3.985000 ;
      RECT 29.241000   3.985000 31.025000   4.055000 ;
      RECT 29.311000   4.055000 31.025000   4.125000 ;
      RECT 29.381000   4.125000 31.025000   4.195000 ;
      RECT 29.451000   4.195000 31.025000   4.265000 ;
      RECT 29.491000   4.503000 31.284000   4.622000 ;
      RECT 29.521000   4.265000 31.025000   4.335000 ;
      RECT 29.591000   4.335000 31.025000   4.405000 ;
      RECT 29.610000   4.622000 31.550000   4.888000 ;
      RECT 29.610000   4.888000 31.550000   6.920000 ;
      RECT 29.661000   4.405000 31.025000   4.475000 ;
      RECT 29.731000   4.475000 31.025000   4.545000 ;
      RECT 29.746000   4.545000 31.025000   4.560000 ;
      RECT 29.750000   4.564000 31.028000   4.635000 ;
      RECT 29.750000   4.635000 31.099000   4.705000 ;
      RECT 29.750000   4.705000 31.169000   4.775000 ;
      RECT 29.750000   4.775000 31.239000   4.845000 ;
      RECT 29.750000   4.845000 31.309000   4.915000 ;
      RECT 29.750000   4.915000 31.379000   4.945000 ;
      RECT 29.750000   4.946000 31.410000   7.060000 ;
      RECT 29.751000   4.561000 31.025000   4.565000 ;
      RECT 29.896000  52.445000 75.950000  52.490000 ;
      RECT 29.896000  52.445000 75.950000  52.490000 ;
      RECT 29.966000  52.375000 75.950000  52.445000 ;
      RECT 29.966000  52.375000 75.950000  52.445000 ;
      RECT 30.036000  52.305000 75.950000  52.375000 ;
      RECT 30.036000  52.305000 75.950000  52.375000 ;
      RECT 30.106000  52.235000 75.950000  52.305000 ;
      RECT 30.106000  52.235000 75.950000  52.305000 ;
      RECT 30.176000  52.165000 75.950000  52.235000 ;
      RECT 30.176000  52.165000 75.950000  52.235000 ;
      RECT 30.246000  52.095000 75.950000  52.165000 ;
      RECT 30.246000  52.095000 75.950000  52.165000 ;
      RECT 30.316000  52.025000 75.950000  52.095000 ;
      RECT 30.316000  52.025000 75.950000  52.095000 ;
      RECT 30.386000  51.955000 75.950000  52.025000 ;
      RECT 30.386000  51.955000 75.950000  52.025000 ;
      RECT 30.456000  51.885000 75.950000  51.955000 ;
      RECT 30.456000  51.885000 75.950000  51.955000 ;
      RECT 30.525000  17.798000 79.180000  36.287000 ;
      RECT 30.525000  36.287000 79.180000  36.552000 ;
      RECT 30.525000  38.178000 79.180000  47.612000 ;
      RECT 30.525000  47.612000 76.090000  50.702000 ;
      RECT 30.525000  50.702000 76.090000  51.618000 ;
      RECT 30.525000  51.618000 76.090000  52.350000 ;
      RECT 30.526000  51.815000 75.950000  51.885000 ;
      RECT 30.526000  51.815000 75.950000  51.885000 ;
      RECT 30.596000  51.745000 75.950000  51.815000 ;
      RECT 30.596000  51.745000 75.950000  51.815000 ;
      RECT 30.665000  17.856000 79.175000  36.229000 ;
      RECT 30.665000  38.236000 79.175000  42.955000 ;
      RECT 30.665000  42.955000 75.950000  52.490000 ;
      RECT 30.665000  42.955000 79.040000  47.554000 ;
      RECT 30.665000  47.554000 75.950000  52.490000 ;
      RECT 30.665000  47.554000 78.969000  47.625000 ;
      RECT 30.665000  47.554000 78.969000  47.625000 ;
      RECT 30.665000  47.625000 78.899000  47.695000 ;
      RECT 30.665000  47.625000 78.899000  47.695000 ;
      RECT 30.665000  47.695000 78.829000  47.765000 ;
      RECT 30.665000  47.695000 78.829000  47.765000 ;
      RECT 30.665000  47.765000 78.759000  47.835000 ;
      RECT 30.665000  47.765000 78.759000  47.835000 ;
      RECT 30.665000  47.835000 78.689000  47.905000 ;
      RECT 30.665000  47.835000 78.689000  47.905000 ;
      RECT 30.665000  47.905000 78.619000  47.975000 ;
      RECT 30.665000  47.905000 78.619000  47.975000 ;
      RECT 30.665000  47.975000 78.549000  48.045000 ;
      RECT 30.665000  47.975000 78.549000  48.045000 ;
      RECT 30.665000  48.045000 78.479000  48.115000 ;
      RECT 30.665000  48.045000 78.479000  48.115000 ;
      RECT 30.665000  48.115000 78.409000  48.185000 ;
      RECT 30.665000  48.115000 78.409000  48.185000 ;
      RECT 30.665000  48.185000 78.339000  48.255000 ;
      RECT 30.665000  48.185000 78.339000  48.255000 ;
      RECT 30.665000  48.255000 78.269000  48.325000 ;
      RECT 30.665000  48.255000 78.269000  48.325000 ;
      RECT 30.665000  48.325000 78.199000  48.395000 ;
      RECT 30.665000  48.325000 78.199000  48.395000 ;
      RECT 30.665000  48.395000 78.129000  48.465000 ;
      RECT 30.665000  48.395000 78.129000  48.465000 ;
      RECT 30.665000  48.465000 78.059000  48.535000 ;
      RECT 30.665000  48.465000 78.059000  48.535000 ;
      RECT 30.665000  48.535000 77.989000  48.605000 ;
      RECT 30.665000  48.535000 77.989000  48.605000 ;
      RECT 30.665000  48.605000 77.919000  48.675000 ;
      RECT 30.665000  48.605000 77.919000  48.675000 ;
      RECT 30.665000  48.675000 77.849000  48.745000 ;
      RECT 30.665000  48.675000 77.849000  48.745000 ;
      RECT 30.665000  48.745000 77.779000  48.815000 ;
      RECT 30.665000  48.745000 77.779000  48.815000 ;
      RECT 30.665000  48.815000 77.709000  48.885000 ;
      RECT 30.665000  48.815000 77.709000  48.885000 ;
      RECT 30.665000  48.885000 77.639000  48.955000 ;
      RECT 30.665000  48.885000 77.639000  48.955000 ;
      RECT 30.665000  48.955000 77.569000  49.025000 ;
      RECT 30.665000  48.955000 77.569000  49.025000 ;
      RECT 30.665000  49.025000 77.499000  49.095000 ;
      RECT 30.665000  49.025000 77.499000  49.095000 ;
      RECT 30.665000  49.095000 77.429000  49.165000 ;
      RECT 30.665000  49.095000 77.429000  49.165000 ;
      RECT 30.665000  49.165000 77.359000  49.235000 ;
      RECT 30.665000  49.165000 77.359000  49.235000 ;
      RECT 30.665000  49.235000 77.289000  49.305000 ;
      RECT 30.665000  49.235000 77.289000  49.305000 ;
      RECT 30.665000  49.305000 77.219000  49.375000 ;
      RECT 30.665000  49.305000 77.219000  49.375000 ;
      RECT 30.665000  49.375000 77.149000  49.445000 ;
      RECT 30.665000  49.375000 77.149000  49.445000 ;
      RECT 30.665000  49.445000 77.079000  49.515000 ;
      RECT 30.665000  49.445000 77.079000  49.515000 ;
      RECT 30.665000  49.515000 77.009000  49.585000 ;
      RECT 30.665000  49.515000 77.009000  49.585000 ;
      RECT 30.665000  49.585000 76.939000  49.655000 ;
      RECT 30.665000  49.585000 76.939000  49.655000 ;
      RECT 30.665000  49.655000 76.869000  49.725000 ;
      RECT 30.665000  49.655000 76.869000  49.725000 ;
      RECT 30.665000  49.725000 76.799000  49.795000 ;
      RECT 30.665000  49.725000 76.799000  49.795000 ;
      RECT 30.665000  49.795000 76.729000  49.865000 ;
      RECT 30.665000  49.795000 76.729000  49.865000 ;
      RECT 30.665000  49.865000 76.659000  49.935000 ;
      RECT 30.665000  49.865000 76.659000  49.935000 ;
      RECT 30.665000  49.935000 76.589000  50.005000 ;
      RECT 30.665000  49.935000 76.589000  50.005000 ;
      RECT 30.665000  50.005000 76.519000  50.075000 ;
      RECT 30.665000  50.005000 76.519000  50.075000 ;
      RECT 30.665000  50.075000 76.449000  50.145000 ;
      RECT 30.665000  50.075000 76.449000  50.145000 ;
      RECT 30.665000  50.145000 76.379000  50.215000 ;
      RECT 30.665000  50.145000 76.379000  50.215000 ;
      RECT 30.665000  50.215000 76.309000  50.285000 ;
      RECT 30.665000  50.215000 76.309000  50.285000 ;
      RECT 30.665000  50.285000 76.239000  50.355000 ;
      RECT 30.665000  50.285000 76.239000  50.355000 ;
      RECT 30.665000  50.355000 76.169000  50.425000 ;
      RECT 30.665000  50.355000 76.169000  50.425000 ;
      RECT 30.665000  50.425000 76.099000  50.495000 ;
      RECT 30.665000  50.425000 76.099000  50.495000 ;
      RECT 30.665000  50.495000 76.029000  50.565000 ;
      RECT 30.665000  50.495000 76.029000  50.565000 ;
      RECT 30.665000  50.565000 75.959000  50.635000 ;
      RECT 30.665000  50.565000 75.959000  50.635000 ;
      RECT 30.665000  50.635000 75.949000  50.645000 ;
      RECT 30.665000  50.635000 75.949000  50.645000 ;
      RECT 30.665000  50.644000 75.950000  51.676000 ;
      RECT 30.665000  51.676000 75.950000  51.745000 ;
      RECT 30.665000  51.676000 75.950000  51.745000 ;
      RECT 30.716000  17.805000 79.175000  17.855000 ;
      RECT 30.716000  17.805000 79.175000  17.855000 ;
      RECT 30.721000  38.180000 79.175000  38.235000 ;
      RECT 30.721000  38.180000 79.175000  38.235000 ;
      RECT 30.736000  36.229000 79.175000  36.300000 ;
      RECT 30.736000  36.229000 79.175000  36.300000 ;
      RECT 30.786000  17.735000 79.175000  17.805000 ;
      RECT 30.786000  17.735000 79.175000  17.805000 ;
      RECT 30.790000  36.552000 79.180000  37.913000 ;
      RECT 30.790000  37.913000 79.180000  38.178000 ;
      RECT 30.791000  38.110000 79.175000  38.180000 ;
      RECT 30.791000  38.110000 79.175000  38.180000 ;
      RECT 30.806000  36.300000 79.175000  36.370000 ;
      RECT 30.806000  36.300000 79.175000  36.370000 ;
      RECT 30.856000  17.665000 79.175000  17.735000 ;
      RECT 30.856000  17.665000 79.175000  17.735000 ;
      RECT 30.861000  38.040000 79.175000  38.110000 ;
      RECT 30.861000  38.040000 79.175000  38.110000 ;
      RECT 30.876000  36.370000 79.175000  36.440000 ;
      RECT 30.876000  36.370000 79.175000  36.440000 ;
      RECT 30.926000  17.595000 79.175000  17.665000 ;
      RECT 30.926000  17.595000 79.175000  17.665000 ;
      RECT 30.930000  17.856000 79.175000  42.955000 ;
      RECT 30.930000  37.971000 79.175000  38.040000 ;
      RECT 30.930000  37.971000 79.175000  38.040000 ;
      RECT 30.931000  36.440000 79.175000  36.495000 ;
      RECT 30.931000  36.440000 79.175000  36.495000 ;
      RECT 30.996000  17.525000 79.175000  17.595000 ;
      RECT 30.996000  17.525000 79.175000  17.595000 ;
      RECT 31.066000  17.455000 79.175000  17.525000 ;
      RECT 31.066000  17.455000 79.175000  17.525000 ;
      RECT 31.136000  17.385000 79.175000  17.455000 ;
      RECT 31.136000  17.385000 79.175000  17.455000 ;
      RECT 31.150000   0.000000 31.675000   2.097000 ;
      RECT 31.150000   2.097000 31.675000   2.622000 ;
      RECT 31.206000  17.315000 79.175000  17.385000 ;
      RECT 31.206000  17.315000 79.175000  17.385000 ;
      RECT 31.211000  17.310000 79.170000  17.315000 ;
      RECT 31.211000  17.310000 79.170000  17.315000 ;
      RECT 31.235000  17.088000 79.180000  17.798000 ;
      RECT 31.276000  17.245000 79.105000  17.310000 ;
      RECT 31.276000  17.245000 79.105000  17.310000 ;
      RECT 31.290000   0.000000 31.535000   2.039000 ;
      RECT 31.341000  17.180000 79.040000  17.245000 ;
      RECT 31.341000  17.180000 79.040000  17.245000 ;
      RECT 31.356000  17.165000 79.040000  17.180000 ;
      RECT 31.356000  17.165000 79.040000  17.180000 ;
      RECT 31.361000   2.039000 31.535000   2.110000 ;
      RECT 31.375000  17.146000 79.040000  17.165000 ;
      RECT 31.375000  17.146000 79.040000  17.165000 ;
      RECT 31.431000   2.110000 31.535000   2.180000 ;
      RECT 31.436000  17.085000 78.979000  17.145000 ;
      RECT 31.436000  17.085000 78.979000  17.145000 ;
      RECT 31.501000   2.180000 31.535000   2.250000 ;
      RECT 31.506000  17.015000 78.909000  17.085000 ;
      RECT 31.506000  17.015000 78.909000  17.085000 ;
      RECT 31.576000  16.945000 78.839000  17.015000 ;
      RECT 31.576000  16.945000 78.839000  17.015000 ;
      RECT 31.646000  16.875000 78.769000  16.945000 ;
      RECT 31.646000  16.875000 78.769000  16.945000 ;
      RECT 31.705000   4.105000 45.105000   4.277000 ;
      RECT 31.705000   4.277000 45.105000   4.662000 ;
      RECT 31.716000  16.805000 78.699000  16.875000 ;
      RECT 31.716000  16.805000 78.699000  16.875000 ;
      RECT 31.786000  16.735000 78.629000  16.805000 ;
      RECT 31.786000  16.735000 78.629000  16.805000 ;
      RECT 31.856000  16.665000 78.559000  16.735000 ;
      RECT 31.856000  16.665000 78.559000  16.735000 ;
      RECT 31.926000  16.595000 78.489000  16.665000 ;
      RECT 31.926000  16.595000 78.489000  16.665000 ;
      RECT 31.940000  16.383000 79.180000  17.088000 ;
      RECT 31.941000   4.245000 44.965000   4.315000 ;
      RECT 31.995000  16.526000 78.420000  16.595000 ;
      RECT 31.995000  16.526000 78.420000  16.595000 ;
      RECT 32.011000   4.315000 44.965000   4.385000 ;
      RECT 32.021000  16.500000 78.420000  16.525000 ;
      RECT 32.021000  16.500000 78.420000  16.525000 ;
      RECT 32.081000   4.385000 44.965000   4.455000 ;
      RECT 32.090000   4.662000 45.105000   5.148000 ;
      RECT 32.090000   5.148000 45.715000   5.758000 ;
      RECT 32.090000   5.758000 45.715000   6.920000 ;
      RECT 32.090000   6.920000 78.570000  10.112000 ;
      RECT 32.090000  10.112000 78.475000  10.207000 ;
      RECT 32.090000  10.207000 78.475000  16.233000 ;
      RECT 32.090000  16.233000 78.475000  16.383000 ;
      RECT 32.091000  16.430000 78.420000  16.500000 ;
      RECT 32.091000  16.430000 78.420000  16.500000 ;
      RECT 32.151000   4.455000 44.965000   4.525000 ;
      RECT 32.161000  16.360000 78.420000  16.430000 ;
      RECT 32.161000  16.360000 78.420000  16.430000 ;
      RECT 32.215000   0.000000 35.320000   1.842000 ;
      RECT 32.215000   1.842000 34.995000   2.167000 ;
      RECT 32.215000   2.167000 34.995000   4.025000 ;
      RECT 32.215000   4.025000 45.105000   4.105000 ;
      RECT 32.221000   4.525000 44.965000   4.595000 ;
      RECT 32.230000   4.245000 44.965000   4.604000 ;
      RECT 32.230000   4.604000 44.965000   5.206000 ;
      RECT 32.230000   5.206000 44.965000   5.275000 ;
      RECT 32.230000   5.206000 44.965000   5.275000 ;
      RECT 32.230000   5.275000 45.034000   5.345000 ;
      RECT 32.230000   5.275000 45.034000   5.345000 ;
      RECT 32.230000   5.345000 45.104000   5.415000 ;
      RECT 32.230000   5.345000 45.104000   5.415000 ;
      RECT 32.230000   5.415000 45.174000   5.485000 ;
      RECT 32.230000   5.415000 45.174000   5.485000 ;
      RECT 32.230000   5.485000 45.244000   5.555000 ;
      RECT 32.230000   5.485000 45.244000   5.555000 ;
      RECT 32.230000   5.555000 45.314000   5.625000 ;
      RECT 32.230000   5.555000 45.314000   5.625000 ;
      RECT 32.230000   5.625000 45.384000   5.695000 ;
      RECT 32.230000   5.625000 45.384000   5.695000 ;
      RECT 32.230000   5.695000 45.454000   5.765000 ;
      RECT 32.230000   5.695000 45.454000   5.765000 ;
      RECT 32.230000   5.765000 45.524000   5.815000 ;
      RECT 32.230000   5.765000 45.524000   5.815000 ;
      RECT 32.230000   5.816000 45.575000   7.060000 ;
      RECT 32.230000   7.060000 78.420000  16.291000 ;
      RECT 32.230000   7.060000 78.420000  16.291000 ;
      RECT 32.230000   7.060000 78.420000  16.291000 ;
      RECT 32.230000   7.060000 78.420000  16.291000 ;
      RECT 32.230000   7.060000 78.420000  16.291000 ;
      RECT 32.230000   7.060000 78.430000   8.230000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.365000 78.565000   9.910000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.045000 78.430000  10.054000 ;
      RECT 32.230000  10.054000 78.424000  10.060000 ;
      RECT 32.230000  10.054000 78.424000  10.060000 ;
      RECT 32.230000  10.060000 78.419000  10.065000 ;
      RECT 32.230000  10.060000 78.419000  10.065000 ;
      RECT 32.230000  10.064000 78.420000  16.291000 ;
      RECT 32.230000  10.064000 78.420000  17.856000 ;
      RECT 32.230000  16.291000 78.420000  16.360000 ;
      RECT 32.230000  16.291000 78.420000  16.360000 ;
      RECT 32.231000   4.595000 44.965000   4.605000 ;
      RECT 32.355000   0.000000 35.180000   1.784000 ;
      RECT 32.355000   1.784000 35.109000   1.855000 ;
      RECT 32.355000   1.855000 35.039000   1.925000 ;
      RECT 32.355000   1.925000 34.969000   1.995000 ;
      RECT 32.355000   1.995000 34.899000   2.065000 ;
      RECT 32.355000   2.065000 34.854000   2.110000 ;
      RECT 32.355000   2.109000 34.855000   4.165000 ;
      RECT 32.355000   4.165000 44.965000   4.245000 ;
      RECT 35.535000   2.393000 38.250000   3.855000 ;
      RECT 35.535000   3.855000 45.105000   4.025000 ;
      RECT 35.675000   2.451000 38.110000   3.995000 ;
      RECT 35.675000   3.995000 44.965000   4.165000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.721000   2.405000 38.110000   2.450000 ;
      RECT 35.791000   2.335000 38.110000   2.405000 ;
      RECT 35.860000   0.000000 38.250000   2.068000 ;
      RECT 35.860000   2.068000 38.250000   2.393000 ;
      RECT 35.861000   2.265000 38.110000   2.335000 ;
      RECT 35.931000   2.195000 38.110000   2.265000 ;
      RECT 36.000000   0.000000 38.110000   2.126000 ;
      RECT 36.000000   2.126000 38.110000   2.195000 ;
      RECT 38.790000   0.000000 45.105000   3.855000 ;
      RECT 38.930000   0.000000 44.965000   3.995000 ;
      RECT 38.930000   0.000000 44.965000   4.604000 ;
      RECT 38.930000   0.000000 44.965000   5.206000 ;
      RECT 38.930000   0.000000 44.965000   5.206000 ;
      RECT 38.930000   0.000000 44.965000   5.206000 ;
      RECT 38.930000   0.000000 44.965000   5.206000 ;
      RECT 38.930000   0.000000 44.965000   5.206000 ;
      RECT 38.930000   0.000000 44.965000   5.206000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 45.645000   0.000000 49.715000   0.222000 ;
      RECT 45.645000   0.222000 49.450000   0.487000 ;
      RECT 45.645000   0.487000 49.450000   0.965000 ;
      RECT 45.645000   0.965000 66.400000   1.137000 ;
      RECT 45.645000   1.137000 66.400000   1.615000 ;
      RECT 45.645000   1.615000 68.135000   4.100000 ;
      RECT 45.645000   4.100000 77.010000   4.922000 ;
      RECT 45.645000   4.922000 77.010000   5.375000 ;
      RECT 45.785000   0.000000 49.310000   0.164000 ;
      RECT 45.785000   0.164000 49.310000   0.429000 ;
      RECT 45.785000   0.164000 49.504000   0.235000 ;
      RECT 45.785000   0.235000 49.434000   0.305000 ;
      RECT 45.785000   0.305000 49.364000   0.375000 ;
      RECT 45.785000   0.375000 49.309000   0.430000 ;
      RECT 45.785000   0.429000 49.310000   1.105000 ;
      RECT 45.785000   1.105000 66.260000   4.864000 ;
      RECT 45.785000   1.105000 66.260000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.240000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   1.755000 67.995000   4.864000 ;
      RECT 45.785000   4.240000 76.870000   4.864000 ;
      RECT 45.856000   4.864000 76.870000   4.935000 ;
      RECT 45.856000   4.864000 76.870000   4.935000 ;
      RECT 45.926000   4.935000 76.870000   5.005000 ;
      RECT 45.926000   4.935000 76.870000   5.005000 ;
      RECT 45.996000   5.005000 76.870000   5.075000 ;
      RECT 45.996000   5.005000 76.870000   5.075000 ;
      RECT 46.066000   5.075000 76.870000   5.145000 ;
      RECT 46.066000   5.075000 76.870000   5.145000 ;
      RECT 46.098000   5.375000 78.570000   5.532000 ;
      RECT 46.136000   5.145000 76.870000   5.215000 ;
      RECT 46.136000   5.145000 76.870000   5.215000 ;
      RECT 46.206000   5.215000 76.870000   5.285000 ;
      RECT 46.206000   5.215000 76.870000   5.285000 ;
      RECT 46.255000   5.532000 78.570000   6.920000 ;
      RECT 46.276000   5.285000 76.870000   5.355000 ;
      RECT 46.276000   5.285000 76.870000   5.355000 ;
      RECT 46.346000   5.355000 76.870000   5.425000 ;
      RECT 46.346000   5.355000 76.870000   5.425000 ;
      RECT 46.395000   5.474000 76.870000   5.515000 ;
      RECT 46.395000   5.515000 78.430000   7.060000 ;
      RECT 46.396000   5.425000 76.870000   5.475000 ;
      RECT 46.396000   5.425000 76.870000   5.475000 ;
      RECT 49.310000   0.000000 49.575000   0.164000 ;
      RECT 50.255000   0.000000 66.695000   0.242000 ;
      RECT 50.255000   0.242000 66.695000   0.487000 ;
      RECT 50.395000   0.000000 50.640000   0.184000 ;
      RECT 50.466000   0.184000 66.555000   0.255000 ;
      RECT 50.500000   0.487000 66.695000   0.842000 ;
      RECT 50.500000   0.842000 66.572000   0.965000 ;
      RECT 50.536000   0.255000 66.555000   0.325000 ;
      RECT 50.606000   0.325000 66.555000   0.395000 ;
      RECT 50.640000   0.000000 66.260000   4.864000 ;
      RECT 50.640000   0.784000 66.484000   0.855000 ;
      RECT 50.640000   0.855000 66.414000   0.925000 ;
      RECT 50.640000   0.925000 66.344000   0.995000 ;
      RECT 50.640000   0.995000 66.274000   1.065000 ;
      RECT 50.640000   1.065000 66.259000   1.080000 ;
      RECT 50.641000   0.395000 66.555000   0.430000 ;
      RECT 66.260000   0.000000 66.555000   0.184000 ;
      RECT 66.260000   0.429000 66.555000   0.784000 ;
      RECT 67.235000   0.000000 68.135000   0.872000 ;
      RECT 67.235000   0.872000 68.135000   1.137000 ;
      RECT 67.375000   0.000000 67.995000   0.814000 ;
      RECT 67.446000   0.814000 67.995000   0.885000 ;
      RECT 67.500000   1.137000 68.135000   1.615000 ;
      RECT 67.516000   0.885000 67.995000   0.955000 ;
      RECT 67.586000   0.955000 67.995000   1.025000 ;
      RECT 67.640000   1.079000 67.995000   1.755000 ;
      RECT 67.641000   1.025000 67.995000   1.080000 ;
      RECT 69.065000   0.000000 76.140000   2.113000 ;
      RECT 69.065000   2.113000 77.010000   2.983000 ;
      RECT 69.065000   2.983000 77.010000   4.100000 ;
      RECT 69.205000   0.000000 76.000000   3.005000 ;
      RECT 69.205000   2.171000 76.000000   2.240000 ;
      RECT 69.205000   2.171000 76.000000   2.240000 ;
      RECT 69.205000   2.240000 76.069000   2.310000 ;
      RECT 69.205000   2.240000 76.069000   2.310000 ;
      RECT 69.205000   2.310000 76.139000   2.380000 ;
      RECT 69.205000   2.310000 76.139000   2.380000 ;
      RECT 69.205000   2.380000 76.209000   2.450000 ;
      RECT 69.205000   2.380000 76.209000   2.450000 ;
      RECT 69.205000   2.450000 76.279000   2.520000 ;
      RECT 69.205000   2.450000 76.279000   2.520000 ;
      RECT 69.205000   2.520000 76.349000   2.590000 ;
      RECT 69.205000   2.520000 76.349000   2.590000 ;
      RECT 69.205000   2.590000 76.419000   2.660000 ;
      RECT 69.205000   2.590000 76.419000   2.660000 ;
      RECT 69.205000   2.660000 76.489000   2.730000 ;
      RECT 69.205000   2.660000 76.489000   2.730000 ;
      RECT 69.205000   2.730000 76.559000   2.800000 ;
      RECT 69.205000   2.730000 76.559000   2.800000 ;
      RECT 69.205000   2.800000 76.629000   2.870000 ;
      RECT 69.205000   2.800000 76.629000   2.870000 ;
      RECT 69.205000   2.870000 76.699000   2.940000 ;
      RECT 69.205000   2.870000 76.699000   2.940000 ;
      RECT 69.205000   2.940000 76.769000   3.010000 ;
      RECT 69.205000   2.940000 76.769000   3.010000 ;
      RECT 69.205000   3.010000 76.839000   3.040000 ;
      RECT 69.205000   3.010000 76.839000   3.040000 ;
      RECT 69.205000   3.041000 76.870000   4.240000 ;
      RECT 76.570000  50.908000 79.435000  52.367000 ;
      RECT 76.570000  52.367000 79.435000  53.052000 ;
      RECT 76.710000  50.966000 79.435000  52.309000 ;
      RECT 76.776000  50.900000 79.435000  50.965000 ;
      RECT 76.781000  52.309000 79.435000  52.380000 ;
      RECT 76.846000  50.830000 79.435000  50.900000 ;
      RECT 76.851000  52.380000 79.435000  52.450000 ;
      RECT 76.916000  50.760000 79.435000  50.830000 ;
      RECT 76.921000  52.450000 79.435000  52.520000 ;
      RECT 76.986000  50.690000 79.435000  50.760000 ;
      RECT 76.991000  52.520000 79.435000  52.590000 ;
      RECT 77.056000  50.620000 79.435000  50.690000 ;
      RECT 77.060000   0.000000 77.470000   0.927000 ;
      RECT 77.060000   0.927000 77.352000   1.045000 ;
      RECT 77.060000   1.045000 77.250000   1.567000 ;
      RECT 77.060000   1.567000 77.250000   1.605000 ;
      RECT 77.061000  52.590000 79.435000  52.660000 ;
      RECT 77.098000   1.605000 78.570000   2.537000 ;
      RECT 77.126000  50.550000 79.435000  50.620000 ;
      RECT 77.131000  52.660000 79.435000  52.730000 ;
      RECT 77.196000  50.480000 79.435000  50.550000 ;
      RECT 77.201000  52.730000 79.435000  52.800000 ;
      RECT 77.255000  53.052000 79.435000  96.137000 ;
      RECT 77.255000  96.137000 79.435000  96.280000 ;
      RECT 77.266000  50.410000 79.435000  50.480000 ;
      RECT 77.271000  52.800000 79.435000  52.870000 ;
      RECT 77.336000  50.340000 79.435000  50.410000 ;
      RECT 77.341000  52.870000 79.435000  52.940000 ;
      RECT 77.395000  52.994000 79.435000  96.079000 ;
      RECT 77.396000  52.940000 79.435000  52.995000 ;
      RECT 77.398000  96.280000 80.000000  96.365000 ;
      RECT 77.406000  50.270000 79.435000  50.340000 ;
      RECT 77.466000  96.079000 79.435000  96.150000 ;
      RECT 77.476000  50.200000 79.435000  50.270000 ;
      RECT 77.506000   1.745000 78.430000   1.815000 ;
      RECT 77.536000  96.150000 79.435000  96.220000 ;
      RECT 77.546000  50.130000 79.435000  50.200000 ;
      RECT 77.576000   1.815000 78.430000   1.885000 ;
      RECT 77.596000  96.220000 79.435000  96.280000 ;
      RECT 77.616000  50.060000 79.435000  50.130000 ;
      RECT 77.646000   1.885000 78.430000   1.955000 ;
      RECT 77.666000  96.280000 80.000000  96.350000 ;
      RECT 77.686000  49.990000 79.435000  50.060000 ;
      RECT 77.716000   1.955000 78.430000   2.025000 ;
      RECT 77.736000  96.350000 80.000000  96.420000 ;
      RECT 77.756000  49.920000 79.435000  49.990000 ;
      RECT 77.786000   2.025000 78.430000   2.095000 ;
      RECT 77.806000  96.420000 80.000000  96.490000 ;
      RECT 77.821000  96.490000 80.000000  96.505000 ;
      RECT 77.826000  49.850000 79.435000  49.920000 ;
      RECT 77.856000   2.095000 78.430000   2.165000 ;
      RECT 77.896000  49.780000 79.435000  49.850000 ;
      RECT 77.926000   2.165000 78.430000   2.235000 ;
      RECT 77.966000  49.710000 79.435000  49.780000 ;
      RECT 77.996000   2.235000 78.430000   2.305000 ;
      RECT 78.010000   0.000000 78.565000   0.817000 ;
      RECT 78.010000   0.817000 78.565000   1.045000 ;
      RECT 78.030000   2.537000 78.570000   5.375000 ;
      RECT 78.036000  49.640000 79.435000  49.710000 ;
      RECT 78.066000   2.305000 78.430000   2.375000 ;
      RECT 78.106000  49.570000 79.435000  49.640000 ;
      RECT 78.136000   2.375000 78.430000   2.445000 ;
      RECT 78.150000   0.000000 78.425000   0.759000 ;
      RECT 78.170000   2.479000 78.430000   5.515000 ;
      RECT 78.171000   2.445000 78.430000   2.480000 ;
      RECT 78.176000  49.500000 79.435000  49.570000 ;
      RECT 78.221000   0.759000 78.425000   0.830000 ;
      RECT 78.246000  49.430000 79.435000  49.500000 ;
      RECT 78.291000   0.830000 78.425000   0.900000 ;
      RECT 78.296000   0.900000 78.425000   0.905000 ;
      RECT 78.316000  49.360000 79.435000  49.430000 ;
      RECT 78.350000   1.045000 78.565000   1.273000 ;
      RECT 78.350000   1.273000 78.570000   1.278000 ;
      RECT 78.350000   1.278000 78.570000   1.605000 ;
      RECT 78.386000  49.290000 79.435000  49.360000 ;
      RECT 78.456000  49.220000 79.435000  49.290000 ;
      RECT 78.526000  49.150000 79.435000  49.220000 ;
      RECT 78.596000  49.080000 79.435000  49.150000 ;
      RECT 78.666000  49.010000 79.435000  49.080000 ;
      RECT 78.736000  48.940000 79.435000  49.010000 ;
      RECT 78.806000  48.870000 79.435000  48.940000 ;
      RECT 78.876000  48.800000 79.435000  48.870000 ;
      RECT 78.945000  10.503000 79.435000  16.187000 ;
      RECT 78.945000  16.187000 79.435000  16.677000 ;
      RECT 78.946000  48.730000 79.435000  48.800000 ;
      RECT 79.016000  48.660000 79.435000  48.730000 ;
      RECT 79.045000   0.000000 79.435000   1.067000 ;
      RECT 79.045000   1.067000 79.435000   1.072000 ;
      RECT 79.050000   1.072000 79.435000  10.398000 ;
      RECT 79.050000  10.398000 79.435000  10.503000 ;
      RECT 79.085000  10.561000 79.435000  16.129000 ;
      RECT 79.086000  48.590000 79.435000  48.660000 ;
      RECT 79.136000  10.510000 79.435000  10.560000 ;
      RECT 79.156000  16.129000 79.435000  16.200000 ;
      RECT 79.156000  48.520000 79.435000  48.590000 ;
      RECT 79.185000   0.000000 79.435000   1.009000 ;
      RECT 79.190000   1.014000 79.435000  10.456000 ;
      RECT 79.190000  10.456000 79.435000  10.510000 ;
      RECT 79.191000   1.009000 79.435000   1.015000 ;
      RECT 79.226000  16.200000 79.435000  16.270000 ;
      RECT 79.226000  48.450000 79.435000  48.520000 ;
      RECT 79.296000  16.270000 79.435000  16.340000 ;
      RECT 79.296000  48.380000 79.435000  48.450000 ;
      RECT 79.366000  16.340000 79.435000  16.410000 ;
      RECT 79.366000  48.310000 79.435000  48.380000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.100000 106.585000 ;
      RECT  0.000000 118.955000  0.100000 178.609000 ;
      RECT  0.000000 178.609000  2.961000 181.470000 ;
      RECT  0.000000 178.800000  0.149000 178.950000 ;
      RECT  0.000000 178.950000  0.299000 179.100000 ;
      RECT  0.000000 179.100000  0.449000 179.250000 ;
      RECT  0.000000 179.250000  0.599000 179.400000 ;
      RECT  0.000000 179.400000  0.749000 179.550000 ;
      RECT  0.000000 179.550000  0.899000 179.700000 ;
      RECT  0.000000 179.700000  1.049000 179.850000 ;
      RECT  0.000000 179.850000  1.199000 180.000000 ;
      RECT  0.000000 180.000000  1.349000 180.150000 ;
      RECT  0.000000 180.150000  1.499000 180.300000 ;
      RECT  0.000000 180.300000  1.649000 180.450000 ;
      RECT  0.000000 180.450000  1.799000 180.600000 ;
      RECT  0.000000 180.600000  1.949000 180.750000 ;
      RECT  0.000000 180.750000  2.099000 180.900000 ;
      RECT  0.000000 180.900000  2.249000 181.050000 ;
      RECT  0.000000 181.050000  2.399000 181.200000 ;
      RECT  0.000000 181.200000  2.549000 181.350000 ;
      RECT  0.000000 181.350000  2.699000 181.500000 ;
      RECT  0.000000 181.470000 80.000000 200.000000 ;
      RECT  0.000000 181.500000  2.849000 181.570000 ;
      RECT  0.000000 181.570000  7.970000 184.572000 ;
      RECT  0.000000 184.572000  7.967000 184.575000 ;
      RECT  0.000000 184.575000  3.005000 196.995000 ;
      RECT  0.000000 196.995000 80.000000 200.000000 ;
      RECT  1.320000   0.000000 45.565000  36.929000 ;
      RECT  1.320000  36.929000 46.276000  37.640000 ;
      RECT  1.320000  37.640000 60.310000  47.660000 ;
      RECT  1.320000  47.660000 61.410000  74.309000 ;
      RECT  1.320000  74.309000 62.736000  75.635000 ;
      RECT  1.320000  75.635000 68.390000  76.344000 ;
      RECT  1.320000  76.344000 68.390000 102.210000 ;
      RECT  1.320000 102.210000 78.280000 106.585000 ;
      RECT  1.320000 118.955000 78.280000 176.780000 ;
      RECT  1.320000 176.780000 80.000000 178.111000 ;
      RECT  1.320000 178.111000 80.000000 180.140000 ;
      RECT  1.415000   0.945000 45.465000   1.675000 ;
      RECT  1.420000   0.000000 45.465000   0.945000 ;
      RECT  1.420000   1.675000 45.465000   3.950000 ;
      RECT  1.420000   3.950000  4.425000  36.971000 ;
      RECT  1.420000  36.971000 45.465000  37.120000 ;
      RECT  1.420000  37.120000 45.614000  37.270000 ;
      RECT  1.420000  37.270000 45.764000  37.420000 ;
      RECT  1.420000  37.420000 45.914000  37.570000 ;
      RECT  1.420000  37.570000 46.064000  37.720000 ;
      RECT  1.420000  37.720000 46.214000  37.740000 ;
      RECT  1.420000  37.740000  4.425000  74.351000 ;
      RECT  1.420000  74.351000 61.310000  74.500000 ;
      RECT  1.420000  74.500000 61.459000  74.650000 ;
      RECT  1.420000  74.650000 61.609000  74.800000 ;
      RECT  1.420000  74.800000 61.759000  74.950000 ;
      RECT  1.420000  74.950000 61.909000  75.100000 ;
      RECT  1.420000  75.100000 62.059000  75.250000 ;
      RECT  1.420000  75.250000 62.209000  75.400000 ;
      RECT  1.420000  75.400000 62.359000  75.550000 ;
      RECT  1.420000  75.550000 62.509000  75.700000 ;
      RECT  1.420000  75.700000 62.659000  75.735000 ;
      RECT  1.420000  75.735000 67.639000  75.885000 ;
      RECT  1.420000  75.885000 67.789000  76.035000 ;
      RECT  1.420000  76.035000 67.939000  76.185000 ;
      RECT  1.420000  76.185000 68.089000  76.335000 ;
      RECT  1.420000  76.335000 68.239000  76.385000 ;
      RECT  1.420000  76.386000 68.290000 106.585000 ;
      RECT  1.420000 118.955000  4.462000 121.960000 ;
      RECT  1.420000 121.960000  4.425000 173.875000 ;
      RECT  1.420000 173.875000  4.477000 176.880000 ;
      RECT  1.420000 176.880000  4.477000 176.960000 ;
      RECT  1.420000 176.960000  4.557000 177.040000 ;
      RECT  1.420000 177.038000  7.970000 178.069000 ;
      RECT  1.441000 178.069000 80.000000 178.090000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 178.109000  7.970000 178.145000 ;
      RECT  1.461000 178.090000 80.000000 178.110000 ;
      RECT  1.646000 178.145000 80.000000 178.295000 ;
      RECT  1.796000 178.295000 80.000000 178.445000 ;
      RECT  1.946000 178.445000 80.000000 178.595000 ;
      RECT  2.000000 106.585000 78.280000 118.955000 ;
      RECT  2.096000 178.595000 80.000000 178.745000 ;
      RECT  2.246000 178.745000 80.000000 178.895000 ;
      RECT  2.396000 178.895000 80.000000 179.045000 ;
      RECT  2.546000 179.045000 80.000000 179.195000 ;
      RECT  2.696000 179.195000 80.000000 179.345000 ;
      RECT  2.846000 179.345000 80.000000 179.495000 ;
      RECT  2.996000 179.495000 80.000000 179.645000 ;
      RECT  3.002000 184.572000 76.998000 196.998000 ;
      RECT  3.146000 179.645000 80.000000 179.795000 ;
      RECT  3.296000 179.795000 80.000000 179.945000 ;
      RECT  3.391000 179.945000 80.000000 180.040000 ;
      RECT  4.422000   3.002000 42.463000  38.215000 ;
      RECT  4.422000  38.215000 42.463000  38.365000 ;
      RECT  4.422000  38.215000 42.463000  38.365000 ;
      RECT  4.422000  38.365000 42.613000  38.515000 ;
      RECT  4.422000  38.365000 42.613000  38.515000 ;
      RECT  4.422000  38.515000 42.763000  38.665000 ;
      RECT  4.422000  38.515000 42.763000  38.665000 ;
      RECT  4.422000  38.665000 42.913000  38.815000 ;
      RECT  4.422000  38.665000 42.913000  38.815000 ;
      RECT  4.422000  38.815000 43.063000  38.965000 ;
      RECT  4.422000  38.815000 43.063000  38.965000 ;
      RECT  4.422000  38.965000 43.213000  39.115000 ;
      RECT  4.422000  38.965000 43.213000  39.115000 ;
      RECT  4.422000  39.115000 43.363000  39.265000 ;
      RECT  4.422000  39.115000 43.363000  39.265000 ;
      RECT  4.422000  39.265000 43.513000  39.415000 ;
      RECT  4.422000  39.265000 43.513000  39.415000 ;
      RECT  4.422000  39.415000 43.663000  39.565000 ;
      RECT  4.422000  39.415000 43.663000  39.565000 ;
      RECT  4.422000  39.565000 43.813000  39.715000 ;
      RECT  4.422000  39.565000 43.813000  39.715000 ;
      RECT  4.422000  39.715000 43.963000  39.865000 ;
      RECT  4.422000  39.715000 43.963000  39.865000 ;
      RECT  4.422000  39.865000 44.113000  40.015000 ;
      RECT  4.422000  39.865000 44.113000  40.015000 ;
      RECT  4.422000  40.015000 44.263000  40.165000 ;
      RECT  4.422000  40.015000 44.263000  40.165000 ;
      RECT  4.422000  40.165000 44.413000  40.315000 ;
      RECT  4.422000  40.165000 44.413000  40.315000 ;
      RECT  4.422000  40.315000 44.563000  40.465000 ;
      RECT  4.422000  40.315000 44.563000  40.465000 ;
      RECT  4.422000  40.465000 44.713000  40.615000 ;
      RECT  4.422000  40.465000 44.713000  40.615000 ;
      RECT  4.422000  40.615000 44.863000  40.740000 ;
      RECT  4.422000  40.615000 44.863000  40.740000 ;
      RECT  4.422000  40.742000 57.208000  50.762000 ;
      RECT  4.422000  50.762000 58.308000  75.595000 ;
      RECT  4.422000  75.595000 58.308000  75.745000 ;
      RECT  4.422000  75.595000 58.308000  75.745000 ;
      RECT  4.422000  75.745000 58.458000  75.895000 ;
      RECT  4.422000  75.745000 58.458000  75.895000 ;
      RECT  4.422000  75.895000 58.608000  76.045000 ;
      RECT  4.422000  75.895000 58.608000  76.045000 ;
      RECT  4.422000  76.045000 58.758000  76.195000 ;
      RECT  4.422000  76.045000 58.758000  76.195000 ;
      RECT  4.422000  76.195000 58.908000  76.345000 ;
      RECT  4.422000  76.195000 58.908000  76.345000 ;
      RECT  4.422000  76.345000 59.058000  76.495000 ;
      RECT  4.422000  76.345000 59.058000  76.495000 ;
      RECT  4.422000  76.495000 59.208000  76.645000 ;
      RECT  4.422000  76.495000 59.208000  76.645000 ;
      RECT  4.422000  76.645000 59.358000  76.795000 ;
      RECT  4.422000  76.645000 59.358000  76.795000 ;
      RECT  4.422000  76.795000 59.508000  76.945000 ;
      RECT  4.422000  76.795000 59.508000  76.945000 ;
      RECT  4.422000  76.945000 59.658000  77.095000 ;
      RECT  4.422000  76.945000 59.658000  77.095000 ;
      RECT  4.422000  77.095000 59.808000  77.245000 ;
      RECT  4.422000  77.095000 59.808000  77.245000 ;
      RECT  4.422000  77.245000 59.958000  77.395000 ;
      RECT  4.422000  77.245000 59.958000  77.395000 ;
      RECT  4.422000  77.395000 60.108000  77.545000 ;
      RECT  4.422000  77.395000 60.108000  77.545000 ;
      RECT  4.422000  77.545000 60.258000  77.695000 ;
      RECT  4.422000  77.545000 60.258000  77.695000 ;
      RECT  4.422000  77.695000 60.408000  77.845000 ;
      RECT  4.422000  77.695000 60.408000  77.845000 ;
      RECT  4.422000  77.845000 60.558000  77.995000 ;
      RECT  4.422000  77.845000 60.558000  77.995000 ;
      RECT  4.422000  77.995000 60.708000  78.145000 ;
      RECT  4.422000  77.995000 60.708000  78.145000 ;
      RECT  4.422000  78.145000 60.858000  78.295000 ;
      RECT  4.422000  78.145000 60.858000  78.295000 ;
      RECT  4.422000  78.295000 61.008000  78.445000 ;
      RECT  4.422000  78.295000 61.008000  78.445000 ;
      RECT  4.422000  78.445000 61.158000  78.595000 ;
      RECT  4.422000  78.445000 61.158000  78.595000 ;
      RECT  4.422000  78.595000 61.308000  78.735000 ;
      RECT  4.422000  78.595000 61.308000  78.735000 ;
      RECT  4.422000  78.737000 65.288000 103.583000 ;
      RECT  4.422000 121.957000 75.178000 176.825000 ;
      RECT  4.462000 103.583000 65.288000 105.312000 ;
      RECT  4.462000 105.312000 75.178000 121.957000 ;
      RECT  4.527000 176.825000 75.178000 176.930000 ;
      RECT  4.527000 176.825000 75.178000 176.930000 ;
      RECT  4.632000 176.930000 75.178000 177.035000 ;
      RECT  4.632000 176.930000 75.178000 177.035000 ;
      RECT  4.637000 177.035000 75.178000 177.040000 ;
      RECT  4.637000 177.035000 75.178000 177.040000 ;
      RECT  4.865000 180.140000 80.000000 181.470000 ;
      RECT  4.965000 178.069000  7.970000 178.109000 ;
      RECT  4.965000 178.145000  7.970000 181.570000 ;
      RECT  7.967000 177.038000 75.178000 179.882000 ;
      RECT  7.967000 179.882000 76.998000 184.572000 ;
      RECT 42.460000   3.950000 45.465000  36.971000 ;
      RECT 42.463000  37.740000 52.002000  40.745000 ;
      RECT 46.495000   0.000000 62.520000   5.431000 ;
      RECT 46.495000   5.431000 61.961000   5.990000 ;
      RECT 46.495000   5.990000 59.300000   7.301000 ;
      RECT 46.495000   7.301000 59.300000  11.059000 ;
      RECT 46.495000  11.059000 61.170000  12.929000 ;
      RECT 46.495000  12.929000 61.170000  18.081000 ;
      RECT 46.495000  18.081000 60.310000  18.941000 ;
      RECT 46.495000  18.941000 60.310000  35.570000 ;
      RECT 46.495000  35.570000 47.660000  36.314000 ;
      RECT 46.495000  36.314000 47.880000  36.534000 ;
      RECT 46.495000  36.534000 47.880000  36.541000 ;
      RECT 46.495000  36.541000 47.880000  36.611000 ;
      RECT 46.565000  36.611000 47.781000  36.710000 ;
      RECT 46.595000   0.000000 62.420000   3.005000 ;
      RECT 46.595000   3.005000 49.600000   5.389000 ;
      RECT 46.595000   5.389000 62.269000   5.540000 ;
      RECT 46.595000   5.540000 62.119000   5.690000 ;
      RECT 46.595000   5.690000 61.969000   5.840000 ;
      RECT 46.595000   5.840000 61.919000   5.890000 ;
      RECT 46.595000   5.890000 60.419000   6.040000 ;
      RECT 46.595000   6.040000 60.269000   6.190000 ;
      RECT 46.595000   6.190000 60.119000   6.340000 ;
      RECT 46.595000   6.340000 59.969000   6.490000 ;
      RECT 46.595000   6.490000 59.819000   6.640000 ;
      RECT 46.595000   6.640000 59.669000   6.790000 ;
      RECT 46.595000   6.790000 59.519000   6.940000 ;
      RECT 46.595000   6.940000 59.369000   7.090000 ;
      RECT 46.595000   7.090000 59.219000   7.240000 ;
      RECT 46.595000   7.240000 59.199000   7.260000 ;
      RECT 46.595000   7.259000 59.200000  35.470000 ;
      RECT 46.595000  11.101000 59.200000  11.250000 ;
      RECT 46.595000  11.250000 59.349000  11.400000 ;
      RECT 46.595000  11.400000 59.499000  11.550000 ;
      RECT 46.595000  11.550000 59.649000  11.700000 ;
      RECT 46.595000  11.700000 59.799000  11.850000 ;
      RECT 46.595000  11.850000 59.949000  12.000000 ;
      RECT 46.595000  12.000000 60.099000  12.150000 ;
      RECT 46.595000  12.150000 60.249000  12.300000 ;
      RECT 46.595000  12.300000 60.399000  12.450000 ;
      RECT 46.595000  12.450000 60.549000  12.600000 ;
      RECT 46.595000  12.600000 60.699000  12.750000 ;
      RECT 46.595000  12.750000 60.849000  12.900000 ;
      RECT 46.595000  12.900000 60.999000  12.970000 ;
      RECT 46.595000  18.039000 60.919000  18.190000 ;
      RECT 46.595000  18.190000 60.769000  18.340000 ;
      RECT 46.595000  18.340000 60.619000  18.490000 ;
      RECT 46.595000  18.490000 60.469000  18.640000 ;
      RECT 46.595000  18.640000 60.319000  18.790000 ;
      RECT 46.595000  18.790000 60.209000  18.900000 ;
      RECT 46.595000  35.470000 47.560000  36.356000 ;
      RECT 46.595000  36.356000 47.560000  36.425000 ;
      RECT 46.595000  36.425000 47.629000  36.495000 ;
      RECT 46.595000  36.495000 47.699000  36.500000 ;
      RECT 46.651000  36.499000 47.703000  36.555000 ;
      RECT 46.706000  36.555000 47.759000  36.610000 ;
      RECT 48.311000  37.640000 60.210000  37.740000 ;
      RECT 48.461000  37.490000 60.210000  37.640000 ;
      RECT 48.611000  37.340000 60.210000  37.490000 ;
      RECT 48.761000  37.190000 60.210000  37.340000 ;
      RECT 48.810000  36.544000 60.310000  36.999000 ;
      RECT 48.810000  36.999000 60.310000  37.640000 ;
      RECT 48.910000  36.586000 52.145000  37.041000 ;
      RECT 48.910000  37.041000 60.210000  37.190000 ;
      RECT 49.026000  36.470000 60.210000  36.585000 ;
      RECT 49.040000  35.570000 60.310000  36.314000 ;
      RECT 49.040000  36.314000 60.310000  36.544000 ;
      RECT 49.140000  35.470000 52.145000  36.586000 ;
      RECT 49.140000  36.356000 60.210000  36.470000 ;
      RECT 49.512000  40.685000 57.208000  40.740000 ;
      RECT 49.512000  40.685000 57.208000  40.740000 ;
      RECT 49.597000   3.002000 59.063000   3.150000 ;
      RECT 49.597000   3.002000 59.063000   3.150000 ;
      RECT 49.597000   3.150000 58.913000   3.300000 ;
      RECT 49.597000   3.150000 58.913000   3.300000 ;
      RECT 49.597000   3.300000 58.763000   3.450000 ;
      RECT 49.597000   3.300000 58.763000   3.450000 ;
      RECT 49.597000   3.450000 58.613000   3.600000 ;
      RECT 49.597000   3.450000 58.613000   3.600000 ;
      RECT 49.597000   3.600000 58.463000   3.750000 ;
      RECT 49.597000   3.600000 58.463000   3.750000 ;
      RECT 49.597000   3.750000 58.313000   3.900000 ;
      RECT 49.597000   3.750000 58.313000   3.900000 ;
      RECT 49.597000   3.900000 58.163000   4.050000 ;
      RECT 49.597000   3.900000 58.163000   4.050000 ;
      RECT 49.597000   4.050000 58.013000   4.200000 ;
      RECT 49.597000   4.050000 58.013000   4.200000 ;
      RECT 49.597000   4.200000 57.863000   4.350000 ;
      RECT 49.597000   4.200000 57.863000   4.350000 ;
      RECT 49.597000   4.350000 57.713000   4.500000 ;
      RECT 49.597000   4.350000 57.713000   4.500000 ;
      RECT 49.597000   4.500000 57.563000   4.650000 ;
      RECT 49.597000   4.500000 57.563000   4.650000 ;
      RECT 49.597000   4.650000 57.413000   4.800000 ;
      RECT 49.597000   4.650000 57.413000   4.800000 ;
      RECT 49.597000   4.800000 57.263000   4.950000 ;
      RECT 49.597000   4.800000 57.263000   4.950000 ;
      RECT 49.597000   4.950000 57.113000   5.100000 ;
      RECT 49.597000   4.950000 57.113000   5.100000 ;
      RECT 49.597000   5.100000 56.963000   5.250000 ;
      RECT 49.597000   5.100000 56.963000   5.250000 ;
      RECT 49.597000   5.250000 56.813000   5.400000 ;
      RECT 49.597000   5.250000 56.813000   5.400000 ;
      RECT 49.597000   5.400000 56.663000   5.550000 ;
      RECT 49.597000   5.400000 56.663000   5.550000 ;
      RECT 49.597000   5.550000 56.513000   5.700000 ;
      RECT 49.597000   5.550000 56.513000   5.700000 ;
      RECT 49.597000   5.700000 56.363000   5.850000 ;
      RECT 49.597000   5.700000 56.363000   5.850000 ;
      RECT 49.597000   5.850000 56.213000   6.000000 ;
      RECT 49.597000   5.850000 56.213000   6.000000 ;
      RECT 49.597000   6.000000 56.198000   6.015000 ;
      RECT 49.597000   6.000000 56.198000   6.015000 ;
      RECT 49.597000   6.015000 56.198000  12.345000 ;
      RECT 49.597000  12.345000 56.198000  12.495000 ;
      RECT 49.597000  12.345000 56.198000  12.495000 ;
      RECT 49.597000  12.495000 56.348000  12.645000 ;
      RECT 49.597000  12.495000 56.348000  12.645000 ;
      RECT 49.597000  12.645000 56.498000  12.795000 ;
      RECT 49.597000  12.645000 56.498000  12.795000 ;
      RECT 49.597000  12.795000 56.648000  12.945000 ;
      RECT 49.597000  12.795000 56.648000  12.945000 ;
      RECT 49.597000  12.945000 56.798000  13.095000 ;
      RECT 49.597000  12.945000 56.798000  13.095000 ;
      RECT 49.597000  13.095000 56.948000  13.245000 ;
      RECT 49.597000  13.095000 56.948000  13.245000 ;
      RECT 49.597000  13.245000 57.098000  13.395000 ;
      RECT 49.597000  13.245000 57.098000  13.395000 ;
      RECT 49.597000  13.395000 57.248000  13.545000 ;
      RECT 49.597000  13.395000 57.248000  13.545000 ;
      RECT 49.597000  13.545000 57.398000  13.695000 ;
      RECT 49.597000  13.545000 57.398000  13.695000 ;
      RECT 49.597000  13.695000 57.548000  13.845000 ;
      RECT 49.597000  13.695000 57.548000  13.845000 ;
      RECT 49.597000  13.845000 57.698000  13.995000 ;
      RECT 49.597000  13.845000 57.698000  13.995000 ;
      RECT 49.597000  13.995000 57.848000  14.145000 ;
      RECT 49.597000  13.995000 57.848000  14.145000 ;
      RECT 49.597000  14.145000 57.998000  14.215000 ;
      RECT 49.597000  14.145000 57.998000  14.215000 ;
      RECT 49.597000  14.215000 58.068000  16.795000 ;
      RECT 49.597000  16.795000 57.918000  16.945000 ;
      RECT 49.597000  16.795000 57.918000  16.945000 ;
      RECT 49.597000  16.945000 57.768000  17.095000 ;
      RECT 49.597000  16.945000 57.768000  17.095000 ;
      RECT 49.597000  17.095000 57.618000  17.245000 ;
      RECT 49.597000  17.095000 57.618000  17.245000 ;
      RECT 49.597000  17.245000 57.468000  17.395000 ;
      RECT 49.597000  17.245000 57.468000  17.395000 ;
      RECT 49.597000  17.395000 57.318000  17.545000 ;
      RECT 49.597000  17.395000 57.318000  17.545000 ;
      RECT 49.597000  17.545000 57.208000  17.655000 ;
      RECT 49.597000  17.545000 57.208000  17.655000 ;
      RECT 49.597000  17.655000 57.208000  32.468000 ;
      RECT 49.662000  40.535000 57.208000  40.685000 ;
      RECT 49.662000  40.535000 57.208000  40.685000 ;
      RECT 49.812000  40.385000 57.208000  40.535000 ;
      RECT 49.812000  40.385000 57.208000  40.535000 ;
      RECT 49.962000  40.235000 57.208000  40.385000 ;
      RECT 49.962000  40.235000 57.208000  40.385000 ;
      RECT 50.112000  40.085000 57.208000  40.235000 ;
      RECT 50.112000  40.085000 57.208000  40.235000 ;
      RECT 50.262000  39.935000 57.208000  40.085000 ;
      RECT 50.262000  39.935000 57.208000  40.085000 ;
      RECT 50.412000  39.785000 57.208000  39.935000 ;
      RECT 50.412000  39.785000 57.208000  39.935000 ;
      RECT 50.562000  39.635000 57.208000  39.785000 ;
      RECT 50.562000  39.635000 57.208000  39.785000 ;
      RECT 50.712000  39.485000 57.208000  39.635000 ;
      RECT 50.712000  39.485000 57.208000  39.635000 ;
      RECT 50.862000  39.335000 57.208000  39.485000 ;
      RECT 50.862000  39.335000 57.208000  39.485000 ;
      RECT 51.012000  39.185000 57.208000  39.335000 ;
      RECT 51.012000  39.185000 57.208000  39.335000 ;
      RECT 51.162000  39.035000 57.208000  39.185000 ;
      RECT 51.162000  39.035000 57.208000  39.185000 ;
      RECT 51.312000  38.885000 57.208000  39.035000 ;
      RECT 51.312000  38.885000 57.208000  39.035000 ;
      RECT 51.462000  38.735000 57.208000  38.885000 ;
      RECT 51.462000  38.735000 57.208000  38.885000 ;
      RECT 51.612000  38.585000 57.208000  38.735000 ;
      RECT 51.612000  38.585000 57.208000  38.735000 ;
      RECT 51.762000  38.435000 57.208000  38.585000 ;
      RECT 51.762000  38.435000 57.208000  38.585000 ;
      RECT 51.912000  37.830000 57.208000  38.285000 ;
      RECT 51.912000  38.285000 57.208000  38.435000 ;
      RECT 51.912000  38.285000 57.208000  38.435000 ;
      RECT 52.027000  37.715000 57.208000  37.830000 ;
      RECT 52.027000  37.715000 57.208000  37.830000 ;
      RECT 52.142000  32.468000 57.208000  37.600000 ;
      RECT 52.142000  37.600000 57.208000  37.715000 ;
      RECT 52.142000  37.600000 57.208000  37.715000 ;
      RECT 56.824000   3.005000 62.420000   5.389000 ;
      RECT 57.205000  18.899000 60.210000  37.041000 ;
      RECT 57.205000  37.740000 60.210000  47.760000 ;
      RECT 57.208000  47.760000 61.310000  50.765000 ;
      RECT 58.065000  12.971000 61.070000  18.039000 ;
      RECT 58.305000  50.765000 61.310000  74.351000 ;
      RECT 60.685000   7.874000 62.520000   7.929000 ;
      RECT 60.685000   7.929000 62.520000  10.486000 ;
      RECT 60.685000  10.486000 62.520000  12.321000 ;
      RECT 60.785000   7.916000 62.365000   7.945000 ;
      RECT 60.785000   7.945000 62.394000   7.970000 ;
      RECT 60.785000   7.971000 62.420000  10.444000 ;
      RECT 60.931000   7.770000 62.219000   7.915000 ;
      RECT 60.936000  10.444000 62.420000  10.595000 ;
      RECT 61.081000   7.620000 62.069000   7.770000 ;
      RECT 61.086000  10.595000 62.420000  10.745000 ;
      RECT 61.189000   7.370000 62.465000   7.874000 ;
      RECT 61.231000   7.470000 61.919000   7.620000 ;
      RECT 61.236000  10.745000 62.420000  10.895000 ;
      RECT 61.386000  10.895000 62.420000  11.045000 ;
      RECT 61.536000  11.045000 62.420000  11.195000 ;
      RECT 61.686000  11.195000 62.420000  11.345000 ;
      RECT 61.695000  19.514000 62.325000  34.721000 ;
      RECT 61.795000  19.556000 62.225000  34.679000 ;
      RECT 61.795000  34.679000 62.074000  34.830000 ;
      RECT 61.795000  34.830000 61.924000  34.980000 ;
      RECT 61.836000  11.345000 62.420000  11.495000 ;
      RECT 61.926000  19.425000 62.225000  19.555000 ;
      RECT 61.986000  11.495000 62.420000  11.645000 ;
      RECT 62.076000  19.275000 62.225000  19.425000 ;
      RECT 62.136000  11.645000 62.420000  11.795000 ;
      RECT 62.286000  11.795000 62.420000  11.945000 ;
      RECT 63.080000  36.324000 78.280000  72.881000 ;
      RECT 63.080000  72.881000 78.280000  73.965000 ;
      RECT 63.180000  36.366000 67.097000  39.371000 ;
      RECT 63.180000  39.371000 66.185000  69.834000 ;
      RECT 63.180000  69.834000 71.941000  72.839000 ;
      RECT 63.196000  36.350000 78.180000  36.365000 ;
      RECT 63.331000  72.839000 78.180000  72.990000 ;
      RECT 63.346000  36.200000 78.180000  36.350000 ;
      RECT 63.481000  72.990000 78.180000  73.140000 ;
      RECT 63.496000  36.050000 78.180000  36.200000 ;
      RECT 63.631000  73.140000 78.180000  73.290000 ;
      RECT 63.646000  35.900000 78.180000  36.050000 ;
      RECT 63.781000  73.290000 78.180000  73.440000 ;
      RECT 63.796000  35.750000 78.180000  35.900000 ;
      RECT 63.931000  73.440000 78.180000  73.590000 ;
      RECT 63.946000  35.600000 78.180000  35.750000 ;
      RECT 63.995000  18.389000 78.280000  35.409000 ;
      RECT 63.995000  35.409000 78.280000  36.324000 ;
      RECT 64.081000  73.590000 78.180000  73.740000 ;
      RECT 64.095000  18.431000 67.292000  21.436000 ;
      RECT 64.095000  21.436000 67.100000  35.451000 ;
      RECT 64.095000  35.451000 78.180000  35.600000 ;
      RECT 64.190000   0.000000 78.280000  18.194000 ;
      RECT 64.190000  18.194000 78.280000  18.389000 ;
      RECT 64.191000  18.335000 78.180000  18.430000 ;
      RECT 64.206000  73.740000 78.180000  73.865000 ;
      RECT 64.290000   0.000000 78.180000   7.455000 ;
      RECT 64.290000   2.690000 78.180000   2.735000 ;
      RECT 64.290000   2.735000 78.225000   2.780000 ;
      RECT 64.290000   2.780000 78.270000   2.785000 ;
      RECT 64.290000   2.785000 78.180000  18.236000 ;
      RECT 64.290000  18.236000 78.180000  18.335000 ;
      RECT 66.182000  37.610000 75.178000  70.863000 ;
      RECT 66.197000  37.595000 75.178000  37.610000 ;
      RECT 66.197000  37.595000 75.178000  37.610000 ;
      RECT 66.347000  37.445000 75.178000  37.595000 ;
      RECT 66.347000  37.445000 75.178000  37.595000 ;
      RECT 66.497000  37.295000 75.178000  37.445000 ;
      RECT 66.497000  37.295000 75.178000  37.445000 ;
      RECT 66.647000  37.145000 75.178000  37.295000 ;
      RECT 66.647000  37.145000 75.178000  37.295000 ;
      RECT 66.797000  36.995000 75.178000  37.145000 ;
      RECT 66.797000  36.995000 75.178000  37.145000 ;
      RECT 66.947000  36.845000 75.178000  36.995000 ;
      RECT 66.947000  36.845000 75.178000  36.995000 ;
      RECT 67.097000  19.675000 75.178000  36.695000 ;
      RECT 67.097000  36.695000 75.178000  36.845000 ;
      RECT 67.097000  36.695000 75.178000  36.845000 ;
      RECT 67.102000  19.670000 75.178000  19.675000 ;
      RECT 67.102000  19.670000 75.178000  19.675000 ;
      RECT 67.197000  19.575000 75.178000  19.670000 ;
      RECT 67.197000  19.575000 75.178000  19.670000 ;
      RECT 67.292000   3.002000 75.178000   3.934000 ;
      RECT 67.292000   3.934000 75.178000   3.980000 ;
      RECT 67.292000   3.934000 75.178000   3.980000 ;
      RECT 67.292000   3.980000 75.224000   4.025000 ;
      RECT 67.292000   3.980000 75.224000   4.025000 ;
      RECT 67.292000   4.025000 75.269000   4.030000 ;
      RECT 67.292000   4.025000 75.269000   4.030000 ;
      RECT 67.292000   4.029000 75.273000   4.453000 ;
      RECT 67.292000   4.453000 75.178000  19.480000 ;
      RECT 67.292000  19.480000 75.178000  19.575000 ;
      RECT 67.292000  19.480000 75.178000  19.575000 ;
      RECT 68.679000  73.965000 78.280000  75.346000 ;
      RECT 68.871000  73.865000 78.180000  74.015000 ;
      RECT 69.021000  74.015000 78.180000  74.165000 ;
      RECT 69.171000  74.165000 78.180000  74.315000 ;
      RECT 69.321000  74.315000 78.180000  74.465000 ;
      RECT 69.471000  74.465000 78.180000  74.615000 ;
      RECT 69.621000  74.615000 78.180000  74.765000 ;
      RECT 69.771000  74.765000 78.180000  74.915000 ;
      RECT 69.921000  74.915000 78.180000  75.065000 ;
      RECT 70.060000  75.346000 78.280000 102.210000 ;
      RECT 70.071000  75.065000 78.180000  75.215000 ;
      RECT 70.112000  70.863000 75.178000  71.010000 ;
      RECT 70.112000  70.863000 75.178000  71.010000 ;
      RECT 70.160000  73.865000 78.180000 118.955000 ;
      RECT 70.161000  75.215000 78.180000  75.305000 ;
      RECT 70.262000  71.010000 75.178000  71.160000 ;
      RECT 70.262000  71.010000 75.178000  71.160000 ;
      RECT 70.412000  71.160000 75.178000  71.310000 ;
      RECT 70.412000  71.160000 75.178000  71.310000 ;
      RECT 70.562000  71.310000 75.178000  71.460000 ;
      RECT 70.562000  71.310000 75.178000  71.460000 ;
      RECT 70.712000  71.460000 75.178000  71.610000 ;
      RECT 70.712000  71.460000 75.178000  71.610000 ;
      RECT 70.862000  71.610000 75.178000  71.760000 ;
      RECT 70.862000  71.610000 75.178000  71.760000 ;
      RECT 71.012000  71.760000 75.178000  71.910000 ;
      RECT 71.012000  71.760000 75.178000  71.910000 ;
      RECT 71.162000  71.910000 75.178000  72.060000 ;
      RECT 71.162000  71.910000 75.178000  72.060000 ;
      RECT 71.312000  72.060000 75.178000  72.210000 ;
      RECT 71.312000  72.060000 75.178000  72.210000 ;
      RECT 71.462000  72.210000 75.178000  72.360000 ;
      RECT 71.462000  72.210000 75.178000  72.360000 ;
      RECT 71.612000  72.360000 75.178000  72.510000 ;
      RECT 71.612000  72.360000 75.178000  72.510000 ;
      RECT 71.762000  72.510000 75.178000  72.660000 ;
      RECT 71.762000  72.510000 75.178000  72.660000 ;
      RECT 71.912000  72.660000 75.178000  72.810000 ;
      RECT 71.912000  72.660000 75.178000  72.810000 ;
      RECT 72.062000  72.810000 75.178000  72.960000 ;
      RECT 72.062000  72.810000 75.178000  72.960000 ;
      RECT 72.212000  72.960000 75.178000  73.110000 ;
      RECT 72.212000  72.960000 75.178000  73.110000 ;
      RECT 72.362000  73.110000 75.178000  73.260000 ;
      RECT 72.362000  73.110000 75.178000  73.260000 ;
      RECT 72.512000  73.260000 75.178000  73.410000 ;
      RECT 72.512000  73.260000 75.178000  73.410000 ;
      RECT 72.662000  73.410000 75.178000  73.560000 ;
      RECT 72.662000  73.410000 75.178000  73.560000 ;
      RECT 72.812000  73.560000 75.178000  73.710000 ;
      RECT 72.812000  73.560000 75.178000  73.710000 ;
      RECT 72.962000  73.710000 75.178000  73.860000 ;
      RECT 72.962000  73.710000 75.178000  73.860000 ;
      RECT 73.112000  73.860000 75.178000  74.010000 ;
      RECT 73.112000  73.860000 75.178000  74.010000 ;
      RECT 73.162000  74.010000 75.178000  74.060000 ;
      RECT 73.162000  74.010000 75.178000  74.060000 ;
      RECT 73.162000  74.060000 75.178000 105.312000 ;
      RECT 75.175000  18.431000 78.180000  35.451000 ;
      RECT 75.175000  36.366000 78.180000  72.839000 ;
      RECT 75.175000 118.955000 78.180000 176.880000 ;
      RECT 75.178000 176.880000 80.000000 179.885000 ;
      RECT 75.270000   2.785000 78.275000   7.455000 ;
      RECT 76.995000 179.885000 80.000000 196.995000 ;
      RECT 78.180000   1.160000 78.190000   1.490000 ;
      RECT 79.870000   0.000000 80.000000 176.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000 80.000000   1.635000 ;
      RECT  0.000000   7.885000  4.675000   8.485000 ;
      RECT  0.000000   7.885000 80.000000   8.485000 ;
      RECT  0.000000  13.935000  4.675000  14.535000 ;
      RECT  0.000000  13.935000 80.000000  14.535000 ;
      RECT  0.000000  18.785000  4.675000  19.385000 ;
      RECT  0.000000  18.785000 80.000000  19.385000 ;
      RECT  0.000000  24.835000  4.675000  25.435000 ;
      RECT  0.000000  24.835000 80.000000  25.435000 ;
      RECT  0.000000  30.885000  4.675000  31.485000 ;
      RECT  0.000000  30.885000 80.000000  31.485000 ;
      RECT  0.000000  35.735000  4.675000  36.335000 ;
      RECT  0.000000  35.735000 80.000000  36.335000 ;
      RECT  0.000000  40.585000  4.675000  41.185000 ;
      RECT  0.000000  40.585000 80.000000  41.185000 ;
      RECT  0.000000  46.635000  4.675000  47.335000 ;
      RECT  0.000000  46.635000 80.000000  47.435000 ;
      RECT  0.000000  57.035000 80.000000  57.835000 ;
      RECT  0.000000  57.135000  4.675000  57.835000 ;
      RECT  0.000000  63.085000  4.675000  63.685000 ;
      RECT  0.000000  63.085000 80.000000  63.685000 ;
      RECT  0.000000  68.935000  4.675000  69.635000 ;
      RECT  0.000000  68.935000 80.000000  69.635000 ;
      RECT  0.000000  95.400000  3.005000 104.215000 ;
      RECT  0.000000  95.400000 80.000000 104.315000 ;
      RECT  0.000000 104.215000  9.484000 104.365000 ;
      RECT  0.000000 104.315000  7.706000 106.285000 ;
      RECT  0.000000 104.365000  9.334000 104.515000 ;
      RECT  0.000000 104.515000  9.184000 104.665000 ;
      RECT  0.000000 104.665000  9.034000 104.815000 ;
      RECT  0.000000 104.815000  8.884000 104.965000 ;
      RECT  0.000000 104.965000  8.734000 105.115000 ;
      RECT  0.000000 105.115000  8.584000 105.265000 ;
      RECT  0.000000 105.265000  8.434000 105.415000 ;
      RECT  0.000000 105.415000  8.284000 105.565000 ;
      RECT  0.000000 105.565000  8.134000 105.715000 ;
      RECT  0.000000 105.715000  7.984000 105.865000 ;
      RECT  0.000000 105.865000  7.834000 106.015000 ;
      RECT  0.000000 106.015000  7.684000 106.165000 ;
      RECT  0.000000 106.165000  7.664000 106.185000 ;
      RECT  0.000000 106.185000  1.600000 106.585000 ;
      RECT  0.000000 106.285000  1.700000 106.585000 ;
      RECT  0.000000 118.955000  1.600000 119.355000 ;
      RECT  0.000000 118.955000  1.700000 119.255000 ;
      RECT  0.000000 119.255000  9.686000 121.550000 ;
      RECT  0.000000 119.355000  7.349000 119.505000 ;
      RECT  0.000000 119.505000  7.499000 119.655000 ;
      RECT  0.000000 119.655000  7.649000 119.805000 ;
      RECT  0.000000 119.805000  7.799000 119.955000 ;
      RECT  0.000000 119.955000  7.949000 120.105000 ;
      RECT  0.000000 120.105000  8.099000 120.255000 ;
      RECT  0.000000 120.255000  8.249000 120.405000 ;
      RECT  0.000000 120.405000  8.399000 120.555000 ;
      RECT  0.000000 120.555000  8.549000 120.705000 ;
      RECT  0.000000 120.705000  8.699000 120.855000 ;
      RECT  0.000000 120.855000  8.849000 121.005000 ;
      RECT  0.000000 121.005000  8.999000 121.155000 ;
      RECT  0.000000 121.155000  9.149000 121.305000 ;
      RECT  0.000000 121.305000  9.299000 121.455000 ;
      RECT  0.000000 121.455000  9.449000 121.605000 ;
      RECT  0.000000 121.550000 80.000000 175.385000 ;
      RECT  0.000000 121.605000  9.599000 121.650000 ;
      RECT  0.000000 121.650000 15.902000 124.655000 ;
      RECT  0.000000 124.655000  3.005000 172.380000 ;
      RECT  0.000000 172.380000  4.672000 175.385000 ;
      RECT  1.365000  14.535000  4.675000  18.785000 ;
      RECT  1.365000  14.535000 78.635000  18.785000 ;
      RECT  1.455000  70.310000  4.675000  94.885000 ;
      RECT  1.570000  47.435000 78.430000  57.035000 ;
      RECT  1.670000   1.635000 78.330000   4.640000 ;
      RECT  1.670000   1.635000 78.330000   7.885000 ;
      RECT  1.670000   4.640000  4.675000   7.885000 ;
      RECT  1.670000   8.485000  4.675000  13.935000 ;
      RECT  1.670000   8.485000 78.330000  13.935000 ;
      RECT  1.670000  19.385000  4.675000  24.835000 ;
      RECT  1.670000  19.385000 78.330000  24.835000 ;
      RECT  1.670000  25.435000  4.675000  30.885000 ;
      RECT  1.670000  25.435000 78.330000  30.885000 ;
      RECT  1.670000  31.485000  4.675000  35.735000 ;
      RECT  1.670000  31.485000 78.330000  35.735000 ;
      RECT  1.670000  36.335000  4.675000  40.585000 ;
      RECT  1.670000  36.335000 78.330000  40.585000 ;
      RECT  1.670000  41.185000  4.675000  46.635000 ;
      RECT  1.670000  41.185000 78.330000  46.635000 ;
      RECT  1.670000  47.335000  4.675000  57.135000 ;
      RECT  1.670000  57.835000  4.675000  63.085000 ;
      RECT  1.670000  57.835000 78.330000  63.085000 ;
      RECT  1.670000  63.685000  4.675000  68.935000 ;
      RECT  1.670000  63.685000 78.330000  68.935000 ;
      RECT  1.670000  69.635000  4.675000  70.310000 ;
      RECT  1.670000  69.635000 78.330000  95.400000 ;
      RECT  1.670000  94.885000 78.330000 104.215000 ;
      RECT  1.670000 175.385000  4.675000 196.995000 ;
      RECT  1.670000 175.385000 78.330000 200.000000 ;
      RECT  1.670000 196.995000 78.330000 200.000000 ;
      RECT  3.002000  98.402000 76.998000 101.213000 ;
      RECT  3.002000 101.213000  8.243000 101.360000 ;
      RECT  3.002000 101.213000  8.243000 101.360000 ;
      RECT  3.002000 101.360000  8.093000 101.510000 ;
      RECT  3.002000 101.360000  8.093000 101.510000 ;
      RECT  3.002000 101.510000  7.943000 101.660000 ;
      RECT  3.002000 101.510000  7.943000 101.660000 ;
      RECT  3.002000 101.660000  7.793000 101.810000 ;
      RECT  3.002000 101.660000  7.793000 101.810000 ;
      RECT  3.002000 101.810000  7.643000 101.960000 ;
      RECT  3.002000 101.810000  7.643000 101.960000 ;
      RECT  3.002000 101.960000  7.493000 102.110000 ;
      RECT  3.002000 101.960000  7.493000 102.110000 ;
      RECT  3.002000 102.110000  7.343000 102.260000 ;
      RECT  3.002000 102.110000  7.343000 102.260000 ;
      RECT  3.002000 102.260000  7.193000 102.410000 ;
      RECT  3.002000 102.260000  7.193000 102.410000 ;
      RECT  3.002000 102.410000  7.043000 102.560000 ;
      RECT  3.002000 102.410000  7.043000 102.560000 ;
      RECT  3.002000 102.560000  6.893000 102.710000 ;
      RECT  3.002000 102.560000  6.893000 102.710000 ;
      RECT  3.002000 102.710000  6.743000 102.860000 ;
      RECT  3.002000 102.710000  6.743000 102.860000 ;
      RECT  3.002000 102.860000  6.593000 103.010000 ;
      RECT  3.002000 102.860000  6.593000 103.010000 ;
      RECT  3.002000 103.010000  6.443000 103.160000 ;
      RECT  3.002000 103.010000  6.443000 103.160000 ;
      RECT  3.002000 103.160000  6.418000 103.185000 ;
      RECT  3.002000 103.160000  6.418000 103.185000 ;
      RECT  3.002000 122.357000  6.105000 122.505000 ;
      RECT  3.002000 122.357000  6.105000 122.505000 ;
      RECT  3.002000 122.505000  6.253000 122.655000 ;
      RECT  3.002000 122.505000  6.253000 122.655000 ;
      RECT  3.002000 122.655000  6.403000 122.805000 ;
      RECT  3.002000 122.655000  6.403000 122.805000 ;
      RECT  3.002000 122.805000  6.553000 122.955000 ;
      RECT  3.002000 122.805000  6.553000 122.955000 ;
      RECT  3.002000 122.955000  6.703000 123.105000 ;
      RECT  3.002000 122.955000  6.703000 123.105000 ;
      RECT  3.002000 123.105000  6.853000 123.255000 ;
      RECT  3.002000 123.105000  6.853000 123.255000 ;
      RECT  3.002000 123.255000  7.003000 123.405000 ;
      RECT  3.002000 123.255000  7.003000 123.405000 ;
      RECT  3.002000 123.405000  7.153000 123.555000 ;
      RECT  3.002000 123.405000  7.153000 123.555000 ;
      RECT  3.002000 123.555000  7.303000 123.705000 ;
      RECT  3.002000 123.555000  7.303000 123.705000 ;
      RECT  3.002000 123.705000  7.453000 123.855000 ;
      RECT  3.002000 123.705000  7.453000 123.855000 ;
      RECT  3.002000 123.855000  7.603000 124.005000 ;
      RECT  3.002000 123.855000  7.603000 124.005000 ;
      RECT  3.002000 124.005000  7.753000 124.155000 ;
      RECT  3.002000 124.005000  7.753000 124.155000 ;
      RECT  3.002000 124.155000  7.903000 124.305000 ;
      RECT  3.002000 124.155000  7.903000 124.305000 ;
      RECT  3.002000 124.305000  8.053000 124.455000 ;
      RECT  3.002000 124.305000  8.053000 124.455000 ;
      RECT  3.002000 124.455000  8.203000 124.605000 ;
      RECT  3.002000 124.455000  8.203000 124.605000 ;
      RECT  3.002000 124.605000  8.353000 124.650000 ;
      RECT  3.002000 124.605000  8.353000 124.650000 ;
      RECT  3.002000 124.652000 76.998000 172.383000 ;
      RECT  4.457000  73.312000 75.328000  91.883000 ;
      RECT  4.672000   3.002000 75.328000  73.312000 ;
      RECT  4.672000  91.883000 75.328000  98.402000 ;
      RECT  4.672000 172.383000 75.328000 196.998000 ;
      RECT  9.880000 121.400000 12.460000 121.650000 ;
      RECT 12.800000 104.315000 80.000000 121.550000 ;
      RECT 12.900000  95.400000 80.000000 121.650000 ;
      RECT 15.902000 101.213000 76.998000 124.652000 ;
      RECT 75.325000   4.640000 78.330000   7.885000 ;
      RECT 75.325000   7.885000 80.000000   8.485000 ;
      RECT 75.325000   8.485000 78.330000  13.935000 ;
      RECT 75.325000  13.935000 80.000000  14.535000 ;
      RECT 75.325000  14.535000 78.635000  18.785000 ;
      RECT 75.325000  18.785000 80.000000  19.385000 ;
      RECT 75.325000  19.385000 78.330000  24.835000 ;
      RECT 75.325000  24.835000 80.000000  25.435000 ;
      RECT 75.325000  25.435000 78.330000  30.885000 ;
      RECT 75.325000  30.885000 80.000000  31.485000 ;
      RECT 75.325000  31.485000 78.330000  35.735000 ;
      RECT 75.325000  35.735000 80.000000  36.335000 ;
      RECT 75.325000  36.335000 78.330000  40.585000 ;
      RECT 75.325000  40.585000 80.000000  41.185000 ;
      RECT 75.325000  41.185000 78.330000  46.635000 ;
      RECT 75.325000  46.635000 80.000000  47.335000 ;
      RECT 75.325000  47.335000 78.330000  57.135000 ;
      RECT 75.325000  57.135000 80.000000  57.835000 ;
      RECT 75.325000  57.835000 78.330000  63.085000 ;
      RECT 75.325000  63.085000 80.000000  63.685000 ;
      RECT 75.325000  63.685000 78.330000  68.935000 ;
      RECT 75.325000  68.935000 80.000000  69.635000 ;
      RECT 75.325000  69.635000 78.330000  94.885000 ;
      RECT 75.325000 175.385000 78.330000 196.995000 ;
      RECT 75.328000 172.380000 80.000000 175.385000 ;
      RECT 76.995000 121.650000 80.000000 172.380000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 124.670000 ;
      RECT  0.000000 124.670000 31.315000 147.815000 ;
      RECT  0.000000 147.815000 80.000000 200.000000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT 54.455000 124.670000 80.000000 147.815000 ;
  END
END sky130_fd_io__top_gpiov2
END LIBRARY
