# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_lvc_b2b
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;

  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 15.375 1.28 17.72 1.345 ;
        RECT 15.31 1.345 17.655 1.41 ;
        RECT 56.055 1.28 56.565 1.35 ;
        RECT 56.125 1.35 56.565 1.42 ;
        RECT 56.155 1.42 56.565 1.45 ;
        RECT 56.155 1.45 56.565 15.815 ;
        RECT 16.445 2.94 17.065 3.01 ;
        RECT 16.515 3.01 17.065 3.08 ;
        RECT 16.585 3.08 17.065 3.15 ;
        RECT 16.655 3.15 17.065 3.22 ;
        RECT 16.655 3.22 17.065 15.26 ;
        RECT 16.655 15.26 17.065 15.33 ;
        RECT 16.585 15.33 17.065 15.4 ;
        RECT 16.515 15.4 17.065 15.47 ;
        RECT 16.445 15.47 17.065 15.54 ;
        RECT 16.375 15.54 17.065 15.61 ;
        RECT 16.305 15.61 17.065 15.665 ;
        RECT 8.355 2.94 9.405 3.01 ;
        RECT 8.355 3.01 9.335 3.08 ;
        RECT 8.355 3.08 9.265 3.15 ;
        RECT 8.355 3.15 9.195 3.22 ;
        RECT 8.355 3.22 9.125 3.29 ;
        RECT 8.355 15.315 9.125 15.385 ;
        RECT 8.355 15.385 9.195 15.455 ;
        RECT 8.355 15.455 9.265 15.525 ;
        RECT 8.355 15.525 9.335 15.595 ;
        RECT 8.355 15.595 9.405 15.665 ;
        RECT 8.355 3.29 9.125 15.315 ;
        RECT 35.995 1.28 37.225 1.35 ;
        RECT 36.065 1.35 37.155 1.42 ;
        RECT 36.135 1.42 37.085 1.49 ;
        RECT 36.165 1.49 37.055 1.52 ;
        RECT 8.355 1.41 17.585 1.48 ;
        RECT 8.355 1.48 17.515 1.55 ;
        RECT 8.355 1.55 17.445 1.62 ;
        RECT 8.355 1.62 17.375 1.69 ;
        RECT 8.355 1.69 17.305 1.76 ;
        RECT 8.355 1.76 17.235 1.83 ;
        RECT 8.355 1.83 17.165 1.9 ;
        RECT 8.355 1.9 17.095 1.97 ;
        RECT 8.355 1.97 17.065 2 ;
        RECT 8.355 15.815 16.995 15.885 ;
        RECT 8.355 15.885 16.925 15.955 ;
        RECT 8.355 15.955 16.855 16.025 ;
        RECT 8.355 16.025 16.785 16.095 ;
        RECT 8.355 16.095 16.715 16.165 ;
        RECT 8.355 16.165 16.645 16.235 ;
        RECT 8.355 16.235 16.575 16.305 ;
        RECT 8.355 16.305 16.505 16.375 ;
        RECT 8.355 16.375 16.435 16.445 ;
        RECT 8.355 16.445 16.365 16.515 ;
        RECT 8.355 16.515 16.295 16.585 ;
        RECT 8.355 16.585 16.225 16.655 ;
        RECT 8.355 16.655 16.155 16.725 ;
        RECT 8.355 16.725 16.105 16.775 ;
        RECT 8.355 15.665 17.065 15.815 ;
        RECT 8.355 16.775 16.105 18.35 ;
        RECT 16.655 0 56.565 0.07 ;
        RECT 16.585 0.07 56.565 0.14 ;
        RECT 16.515 0.14 56.565 0.21 ;
        RECT 16.445 0.21 56.565 0.28 ;
        RECT 16.375 0.28 56.565 0.35 ;
        RECT 16.305 0.35 56.565 0.42 ;
        RECT 16.235 0.42 56.565 0.49 ;
        RECT 16.165 0.49 56.565 0.56 ;
        RECT 16.095 0.56 56.565 0.63 ;
        RECT 16.025 0.63 56.565 0.7 ;
        RECT 15.955 0.7 56.565 0.77 ;
        RECT 15.885 0.77 56.565 0.84 ;
        RECT 15.815 0.84 56.565 0.91 ;
        RECT 15.745 0.91 56.565 0.98 ;
        RECT 15.675 0.98 56.565 1.05 ;
        RECT 15.605 1.05 56.565 1.12 ;
        RECT 15.535 1.12 56.565 1.19 ;
        RECT 15.465 1.19 56.565 1.26 ;
        RECT 15.395 1.26 56.565 1.28 ;
        RECT 36.165 1.52 37.055 15.815 ;
        RECT 8.355 2 17.065 2.94 ;
    END
  END vssd

  PIN bdy2_b2b
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 20.205 1.64 53.535 1.71 ;
        RECT 20.135 1.71 53.535 1.78 ;
        RECT 20.065 1.78 53.535 1.85 ;
        RECT 19.995 1.85 53.535 1.92 ;
        RECT 19.925 1.92 53.535 1.99 ;
        RECT 19.855 1.99 53.535 2.06 ;
        RECT 19.785 2.06 53.535 2.13 ;
        RECT 19.715 2.13 53.535 2.2 ;
        RECT 19.645 2.2 53.535 2.27 ;
        RECT 19.575 2.27 53.535 2.34 ;
        RECT 19.505 2.34 53.535 2.41 ;
        RECT 19.435 2.41 53.535 2.48 ;
        RECT 19.365 2.48 53.535 2.55 ;
        RECT 19.295 2.55 53.535 2.62 ;
        RECT 19.225 2.62 53.535 2.69 ;
        RECT 19.155 2.69 53.535 2.76 ;
        RECT 19.085 2.76 53.535 2.83 ;
        RECT 19.015 2.83 53.535 2.9 ;
        RECT 18.945 2.9 53.535 2.97 ;
        RECT 18.875 2.97 53.535 3.04 ;
        RECT 18.805 3.04 53.535 3.11 ;
        RECT 18.735 3.11 53.535 3.18 ;
        RECT 18.665 3.18 53.535 3.25 ;
        RECT 18.595 3.25 53.535 3.32 ;
        RECT 18.525 3.32 53.535 3.39 ;
        RECT 18.455 3.39 53.535 3.46 ;
        RECT 18.385 3.46 53.535 3.53 ;
        RECT 18.315 3.53 53.535 3.6 ;
        RECT 18.245 3.6 53.535 3.67 ;
        RECT 18.175 3.67 53.535 3.74 ;
        RECT 18.105 3.74 53.535 3.81 ;
        RECT 18.035 3.81 53.535 3.88 ;
        RECT 17.965 3.88 53.535 3.95 ;
        RECT 17.895 3.95 53.535 4.02 ;
        RECT 17.825 4.02 53.535 4.09 ;
        RECT 17.755 4.09 53.535 4.16 ;
        RECT 17.685 4.16 53.535 4.215 ;
        RECT 22.575 0 53.535 0.07 ;
        RECT 22.505 0.07 53.535 0.14 ;
        RECT 22.435 0.14 53.535 0.21 ;
        RECT 22.365 0.21 53.535 0.28 ;
        RECT 22.295 0.28 53.535 0.35 ;
        RECT 22.225 0.35 53.535 0.42 ;
        RECT 22.155 0.42 53.535 0.49 ;
        RECT 22.085 0.49 53.535 0.56 ;
        RECT 22.015 0.56 53.535 0.63 ;
        RECT 21.945 0.63 53.535 0.7 ;
        RECT 21.875 0.7 53.535 0.77 ;
        RECT 21.805 0.77 53.535 0.84 ;
        RECT 21.735 0.84 53.535 0.91 ;
        RECT 21.665 0.91 53.535 0.98 ;
        RECT 21.595 0.98 53.535 1.05 ;
        RECT 21.525 1.05 53.535 1.12 ;
        RECT 21.455 1.12 53.535 1.19 ;
        RECT 21.385 1.19 53.535 1.26 ;
        RECT 21.315 1.26 53.535 1.33 ;
        RECT 21.245 1.33 53.535 1.4 ;
        RECT 21.175 1.4 53.535 1.47 ;
        RECT 21.105 1.47 53.535 1.54 ;
        RECT 21.035 1.54 53.535 1.61 ;
        RECT 20.965 1.61 53.535 1.64 ;
        RECT 17.63 4.215 53.535 8.64 ;
    END
  END bdy2_b2b

  PIN src_bdy_lvc2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 66 74.43 68.01 98.56 ;
        RECT 65.27 73.63 68.74 73.7 ;
        RECT 65.34 73.7 68.67 73.77 ;
        RECT 65.41 73.77 68.6 73.84 ;
        RECT 65.48 73.84 68.53 73.91 ;
        RECT 65.55 73.91 68.46 73.98 ;
        RECT 65.62 73.98 68.39 74.05 ;
        RECT 65.69 74.05 68.32 74.12 ;
        RECT 65.76 74.12 68.25 74.19 ;
        RECT 65.83 74.19 68.18 74.26 ;
        RECT 65.9 74.26 68.11 74.33 ;
        RECT 65.97 74.33 68.04 74.4 ;
        RECT 66 74.4 68.01 74.43 ;
        RECT 16.135 70.99 74.7 73.63 ;
        RECT 65.995 69.94 74.7 70.01 ;
        RECT 65.925 70.01 74.7 70.08 ;
        RECT 65.855 70.08 74.7 70.15 ;
        RECT 65.785 70.15 74.7 70.22 ;
        RECT 65.715 70.22 74.7 70.29 ;
        RECT 65.645 70.29 74.7 70.36 ;
        RECT 65.575 70.36 74.7 70.43 ;
        RECT 65.505 70.43 74.7 70.5 ;
        RECT 65.435 70.5 74.7 70.57 ;
        RECT 65.365 70.57 74.7 70.64 ;
        RECT 65.295 70.64 74.7 70.71 ;
        RECT 65.225 70.71 74.7 70.78 ;
        RECT 65.155 70.78 74.7 70.85 ;
        RECT 65.085 70.85 74.7 70.92 ;
        RECT 65.015 70.92 74.7 70.99 ;
        RECT 65.995 64.68 74.7 69.94 ;
        RECT 65.015 63.63 74.7 63.7 ;
        RECT 65.085 63.7 74.7 63.77 ;
        RECT 65.155 63.77 74.7 63.84 ;
        RECT 65.225 63.84 74.7 63.91 ;
        RECT 65.295 63.91 74.7 63.98 ;
        RECT 65.365 63.98 74.7 64.05 ;
        RECT 65.435 64.05 74.7 64.12 ;
        RECT 65.505 64.12 74.7 64.19 ;
        RECT 65.575 64.19 74.7 64.26 ;
        RECT 65.645 64.26 74.7 64.33 ;
        RECT 65.715 64.33 74.7 64.4 ;
        RECT 65.785 64.4 74.7 64.47 ;
        RECT 65.855 64.47 74.7 64.54 ;
        RECT 65.925 64.54 74.7 64.61 ;
        RECT 65.995 64.61 74.7 64.68 ;
        RECT 16.135 60.99 74.7 63.63 ;
        RECT 65.995 59.94 74.7 60.01 ;
        RECT 65.925 60.01 74.7 60.08 ;
        RECT 65.855 60.08 74.7 60.15 ;
        RECT 65.785 60.15 74.7 60.22 ;
        RECT 65.715 60.22 74.7 60.29 ;
        RECT 65.645 60.29 74.7 60.36 ;
        RECT 65.575 60.36 74.7 60.43 ;
        RECT 65.505 60.43 74.7 60.5 ;
        RECT 65.435 60.5 74.7 60.57 ;
        RECT 65.365 60.57 74.7 60.64 ;
        RECT 65.295 60.64 74.7 60.71 ;
        RECT 65.225 60.71 74.7 60.78 ;
        RECT 65.155 60.78 74.7 60.85 ;
        RECT 65.085 60.85 74.7 60.92 ;
        RECT 65.015 60.92 74.7 60.99 ;
        RECT 65.995 54.685 74.7 59.94 ;
        RECT 65.03 53.65 74.7 53.72 ;
        RECT 65.1 53.72 74.7 53.79 ;
        RECT 65.17 53.79 74.7 53.86 ;
        RECT 65.24 53.86 74.7 53.93 ;
        RECT 65.31 53.93 74.7 54 ;
        RECT 65.38 54 74.7 54.07 ;
        RECT 65.45 54.07 74.7 54.14 ;
        RECT 65.52 54.14 74.7 54.21 ;
        RECT 65.59 54.21 74.7 54.28 ;
        RECT 65.66 54.28 74.7 54.35 ;
        RECT 65.73 54.35 74.7 54.42 ;
        RECT 65.8 54.42 74.7 54.49 ;
        RECT 65.87 54.49 74.7 54.56 ;
        RECT 65.94 54.56 74.7 54.63 ;
        RECT 65.995 54.63 74.7 54.685 ;
        RECT 16.135 51.01 74.7 53.65 ;
        RECT 66 49.955 74.7 50.025 ;
        RECT 65.93 50.025 74.7 50.095 ;
        RECT 65.86 50.095 74.7 50.165 ;
        RECT 65.79 50.165 74.7 50.235 ;
        RECT 65.72 50.235 74.7 50.305 ;
        RECT 65.65 50.305 74.7 50.375 ;
        RECT 65.58 50.375 74.7 50.445 ;
        RECT 65.51 50.445 74.7 50.515 ;
        RECT 65.44 50.515 74.7 50.585 ;
        RECT 65.37 50.585 74.7 50.655 ;
        RECT 65.3 50.655 74.7 50.725 ;
        RECT 65.23 50.725 74.7 50.795 ;
        RECT 65.16 50.795 74.7 50.865 ;
        RECT 65.09 50.865 74.7 50.935 ;
        RECT 65.02 50.935 74.7 51.005 ;
        RECT 64.95 51.005 74.7 51.01 ;
        RECT 66 44.67 74.7 49.955 ;
        RECT 65.03 43.63 74.7 43.7 ;
        RECT 65.1 43.7 74.7 43.77 ;
        RECT 65.17 43.77 74.7 43.84 ;
        RECT 65.24 43.84 74.7 43.91 ;
        RECT 65.31 43.91 74.7 43.98 ;
        RECT 65.38 43.98 74.7 44.05 ;
        RECT 65.45 44.05 74.7 44.12 ;
        RECT 65.52 44.12 74.7 44.19 ;
        RECT 65.59 44.19 74.7 44.26 ;
        RECT 65.66 44.26 74.7 44.33 ;
        RECT 65.73 44.33 74.7 44.4 ;
        RECT 65.8 44.4 74.7 44.47 ;
        RECT 65.87 44.47 74.7 44.54 ;
        RECT 65.94 44.54 74.7 44.61 ;
        RECT 66 44.61 74.7 44.67 ;
        RECT 16.135 40.99 74.7 43.63 ;
        RECT 66 39.935 74.7 40.005 ;
        RECT 65.93 40.005 74.7 40.075 ;
        RECT 65.86 40.075 74.7 40.145 ;
        RECT 65.79 40.145 74.7 40.215 ;
        RECT 65.72 40.215 74.7 40.285 ;
        RECT 65.65 40.285 74.7 40.355 ;
        RECT 65.58 40.355 74.7 40.425 ;
        RECT 65.51 40.425 74.7 40.495 ;
        RECT 65.44 40.495 74.7 40.565 ;
        RECT 65.37 40.565 74.7 40.635 ;
        RECT 65.3 40.635 74.7 40.705 ;
        RECT 65.23 40.705 74.7 40.775 ;
        RECT 65.16 40.775 74.7 40.845 ;
        RECT 65.09 40.845 74.7 40.915 ;
        RECT 65.02 40.915 74.7 40.985 ;
        RECT 64.95 40.985 74.7 40.99 ;
        RECT 66 34.69 74.7 39.935 ;
        RECT 65.03 33.65 74.7 33.72 ;
        RECT 65.1 33.72 74.7 33.79 ;
        RECT 65.17 33.79 74.7 33.86 ;
        RECT 65.24 33.86 74.7 33.93 ;
        RECT 65.31 33.93 74.7 34 ;
        RECT 65.38 34 74.7 34.07 ;
        RECT 65.45 34.07 74.7 34.14 ;
        RECT 65.52 34.14 74.7 34.21 ;
        RECT 65.59 34.21 74.7 34.28 ;
        RECT 65.66 34.28 74.7 34.35 ;
        RECT 65.73 34.35 74.7 34.42 ;
        RECT 65.8 34.42 74.7 34.49 ;
        RECT 65.87 34.49 74.7 34.56 ;
        RECT 65.94 34.56 74.7 34.63 ;
        RECT 66 34.63 74.7 34.69 ;
        RECT 16.135 31.01 74.7 33.65 ;
        RECT 66 29.88 74.7 29.95 ;
        RECT 65.93 29.95 74.7 30.02 ;
        RECT 65.86 30.02 74.7 30.09 ;
        RECT 65.79 30.09 74.7 30.16 ;
        RECT 65.72 30.16 74.7 30.23 ;
        RECT 65.65 30.23 74.7 30.3 ;
        RECT 65.58 30.3 74.7 30.37 ;
        RECT 65.51 30.37 74.7 30.44 ;
        RECT 65.44 30.44 74.7 30.51 ;
        RECT 65.37 30.51 74.7 30.58 ;
        RECT 65.3 30.58 74.7 30.65 ;
        RECT 65.23 30.65 74.7 30.72 ;
        RECT 65.16 30.72 74.7 30.79 ;
        RECT 65.09 30.79 74.7 30.86 ;
        RECT 65.02 30.86 74.7 30.93 ;
        RECT 64.95 30.93 74.7 31 ;
        RECT 64.88 31 74.7 31.01 ;
        RECT 66 25.44 74.7 29.88 ;
        RECT 62.325 21.695 74.7 21.765 ;
        RECT 62.395 21.765 74.7 21.835 ;
        RECT 62.465 21.835 74.7 21.905 ;
        RECT 62.535 21.905 74.7 21.975 ;
        RECT 62.605 21.975 74.7 22.045 ;
        RECT 62.675 22.045 74.7 22.115 ;
        RECT 62.745 22.115 74.7 22.185 ;
        RECT 62.815 22.185 74.7 22.255 ;
        RECT 62.885 22.255 74.7 22.325 ;
        RECT 62.955 22.325 74.7 22.395 ;
        RECT 63.025 22.395 74.7 22.465 ;
        RECT 63.095 22.465 74.7 22.535 ;
        RECT 63.165 22.535 74.7 22.605 ;
        RECT 63.235 22.605 74.7 22.675 ;
        RECT 63.305 22.675 74.7 22.745 ;
        RECT 63.375 22.745 74.7 22.815 ;
        RECT 63.445 22.815 74.7 22.885 ;
        RECT 63.515 22.885 74.7 22.955 ;
        RECT 63.585 22.955 74.7 23.025 ;
        RECT 63.655 23.025 74.7 23.095 ;
        RECT 63.725 23.095 74.7 23.165 ;
        RECT 63.795 23.165 74.7 23.235 ;
        RECT 63.865 23.235 74.7 23.305 ;
        RECT 63.935 23.305 74.7 23.375 ;
        RECT 64.005 23.375 74.7 23.445 ;
        RECT 64.075 23.445 74.7 23.515 ;
        RECT 64.145 23.515 74.7 23.585 ;
        RECT 64.215 23.585 74.7 23.655 ;
        RECT 64.285 23.655 74.7 23.725 ;
        RECT 64.355 23.725 74.7 23.795 ;
        RECT 64.425 23.795 74.7 23.865 ;
        RECT 64.495 23.865 74.7 23.935 ;
        RECT 64.565 23.935 74.7 24.005 ;
        RECT 64.635 24.005 74.7 24.075 ;
        RECT 64.705 24.075 74.7 24.145 ;
        RECT 64.775 24.145 74.7 24.215 ;
        RECT 64.845 24.215 74.7 24.285 ;
        RECT 64.915 24.285 74.7 24.355 ;
        RECT 64.985 24.355 74.7 24.425 ;
        RECT 65.055 24.425 74.7 24.495 ;
        RECT 65.125 24.495 74.7 24.565 ;
        RECT 65.195 24.565 74.7 24.635 ;
        RECT 65.265 24.635 74.7 24.705 ;
        RECT 65.335 24.705 74.7 24.775 ;
        RECT 65.405 24.775 74.7 24.845 ;
        RECT 65.475 24.845 74.7 24.915 ;
        RECT 65.545 24.915 74.7 24.985 ;
        RECT 65.615 24.985 74.7 25.055 ;
        RECT 65.685 25.055 74.7 25.125 ;
        RECT 65.755 25.125 74.7 25.195 ;
        RECT 65.825 25.195 74.7 25.265 ;
        RECT 65.895 25.265 74.7 25.335 ;
        RECT 65.965 25.335 74.7 25.405 ;
        RECT 66 25.405 74.7 25.44 ;
        RECT 54.095 19.99 74.7 21.695 ;
        RECT 56.25 17.835 74.7 17.905 ;
        RECT 56.18 17.905 74.7 17.975 ;
        RECT 56.11 17.975 74.7 18.045 ;
        RECT 56.04 18.045 74.7 18.115 ;
        RECT 55.97 18.115 74.7 18.185 ;
        RECT 55.9 18.185 74.7 18.255 ;
        RECT 55.83 18.255 74.7 18.325 ;
        RECT 55.76 18.325 74.7 18.395 ;
        RECT 55.69 18.395 74.7 18.465 ;
        RECT 55.62 18.465 74.7 18.535 ;
        RECT 55.55 18.535 74.7 18.605 ;
        RECT 55.48 18.605 74.7 18.675 ;
        RECT 55.41 18.675 74.7 18.745 ;
        RECT 55.34 18.745 74.7 18.815 ;
        RECT 55.27 18.815 74.7 18.885 ;
        RECT 55.2 18.885 74.7 18.955 ;
        RECT 55.13 18.955 74.7 19.025 ;
        RECT 55.06 19.025 74.7 19.095 ;
        RECT 54.99 19.095 74.7 19.165 ;
        RECT 54.92 19.165 74.7 19.235 ;
        RECT 54.85 19.235 74.7 19.305 ;
        RECT 54.78 19.305 74.7 19.375 ;
        RECT 54.71 19.375 74.7 19.445 ;
        RECT 54.64 19.445 74.7 19.515 ;
        RECT 54.57 19.515 74.7 19.585 ;
        RECT 54.5 19.585 74.7 19.655 ;
        RECT 54.43 19.655 74.7 19.725 ;
        RECT 54.36 19.725 74.7 19.795 ;
        RECT 54.29 19.795 74.7 19.865 ;
        RECT 54.22 19.865 74.7 19.935 ;
        RECT 54.15 19.935 74.7 19.99 ;
        RECT 56.25 9.04 74.7 17.835 ;
        RECT 54.165 6.885 74.7 6.955 ;
        RECT 54.235 6.955 74.7 7.025 ;
        RECT 54.305 7.025 74.7 7.095 ;
        RECT 54.375 7.095 74.7 7.165 ;
        RECT 54.445 7.165 74.7 7.235 ;
        RECT 54.515 7.235 74.7 7.305 ;
        RECT 54.585 7.305 74.7 7.375 ;
        RECT 54.655 7.375 74.7 7.445 ;
        RECT 54.725 7.445 74.7 7.515 ;
        RECT 54.795 7.515 74.7 7.585 ;
        RECT 54.865 7.585 74.7 7.655 ;
        RECT 54.935 7.655 74.7 7.725 ;
        RECT 55.005 7.725 74.7 7.795 ;
        RECT 55.075 7.795 74.7 7.865 ;
        RECT 55.145 7.865 74.7 7.935 ;
        RECT 55.215 7.935 74.7 8.005 ;
        RECT 55.285 8.005 74.7 8.075 ;
        RECT 55.355 8.075 74.7 8.145 ;
        RECT 55.425 8.145 74.7 8.215 ;
        RECT 55.495 8.215 74.7 8.285 ;
        RECT 55.565 8.285 74.7 8.355 ;
        RECT 55.635 8.355 74.7 8.425 ;
        RECT 55.705 8.425 74.7 8.495 ;
        RECT 55.775 8.495 74.7 8.565 ;
        RECT 55.845 8.565 74.7 8.635 ;
        RECT 55.915 8.635 74.7 8.705 ;
        RECT 55.985 8.705 74.7 8.775 ;
        RECT 56.055 8.775 74.7 8.845 ;
        RECT 56.125 8.845 74.7 8.915 ;
        RECT 56.195 8.915 74.7 8.985 ;
        RECT 56.25 8.985 74.7 9.04 ;
        RECT 54.095 0 74.7 6.885 ;
    END
  END src_bdy_lvc2

  PIN src_bdy_lvc1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.5 190.99 68.01 193.63 ;
        RECT 0.5 189.94 13.96 190.01 ;
        RECT 0.5 190.01 14.03 190.08 ;
        RECT 0.5 190.08 14.1 190.15 ;
        RECT 0.5 190.15 14.17 190.22 ;
        RECT 0.5 190.22 14.24 190.29 ;
        RECT 0.5 190.29 14.31 190.36 ;
        RECT 0.5 190.36 14.38 190.43 ;
        RECT 0.5 190.43 14.45 190.5 ;
        RECT 0.5 190.5 14.52 190.57 ;
        RECT 0.5 190.57 14.59 190.64 ;
        RECT 0.5 190.64 14.66 190.71 ;
        RECT 0.5 190.71 14.73 190.78 ;
        RECT 0.5 190.78 14.8 190.85 ;
        RECT 0.5 190.85 14.87 190.92 ;
        RECT 0.5 190.92 14.94 190.99 ;
        RECT 0.5 184.68 13.96 189.94 ;
        RECT 0.5 183.63 14.94 183.7 ;
        RECT 0.5 183.7 14.87 183.77 ;
        RECT 0.5 183.77 14.8 183.84 ;
        RECT 0.5 183.84 14.73 183.91 ;
        RECT 0.5 183.91 14.66 183.98 ;
        RECT 0.5 183.98 14.59 184.05 ;
        RECT 0.5 184.05 14.52 184.12 ;
        RECT 0.5 184.12 14.45 184.19 ;
        RECT 0.5 184.19 14.38 184.26 ;
        RECT 0.5 184.26 14.31 184.33 ;
        RECT 0.5 184.33 14.24 184.4 ;
        RECT 0.5 184.4 14.17 184.47 ;
        RECT 0.5 184.47 14.1 184.54 ;
        RECT 0.5 184.54 14.03 184.61 ;
        RECT 0.5 184.61 13.96 184.68 ;
        RECT 0.5 180.99 68.01 183.63 ;
        RECT 0.5 179.94 13.96 180.01 ;
        RECT 0.5 180.01 14.03 180.08 ;
        RECT 0.5 180.08 14.1 180.15 ;
        RECT 0.5 180.15 14.17 180.22 ;
        RECT 0.5 180.22 14.24 180.29 ;
        RECT 0.5 180.29 14.31 180.36 ;
        RECT 0.5 180.36 14.38 180.43 ;
        RECT 0.5 180.43 14.45 180.5 ;
        RECT 0.5 180.5 14.52 180.57 ;
        RECT 0.5 180.57 14.59 180.64 ;
        RECT 0.5 180.64 14.66 180.71 ;
        RECT 0.5 180.71 14.73 180.78 ;
        RECT 0.5 180.78 14.8 180.85 ;
        RECT 0.5 180.85 14.87 180.92 ;
        RECT 0.5 180.92 14.94 180.99 ;
        RECT 0.5 174.68 13.96 179.94 ;
        RECT 0.5 173.63 14.94 173.7 ;
        RECT 0.5 173.7 14.87 173.77 ;
        RECT 0.5 173.77 14.8 173.84 ;
        RECT 0.5 173.84 14.73 173.91 ;
        RECT 0.5 173.91 14.66 173.98 ;
        RECT 0.5 173.98 14.59 174.05 ;
        RECT 0.5 174.05 14.52 174.12 ;
        RECT 0.5 174.12 14.45 174.19 ;
        RECT 0.5 174.19 14.38 174.26 ;
        RECT 0.5 174.26 14.31 174.33 ;
        RECT 0.5 174.33 14.24 174.4 ;
        RECT 0.5 174.4 14.17 174.47 ;
        RECT 0.5 174.47 14.1 174.54 ;
        RECT 0.5 174.54 14.03 174.61 ;
        RECT 0.5 174.61 13.96 174.68 ;
        RECT 0.5 170.99 68.01 173.63 ;
        RECT 0.5 169.94 13.96 170.01 ;
        RECT 0.5 170.01 14.03 170.08 ;
        RECT 0.5 170.08 14.1 170.15 ;
        RECT 0.5 170.15 14.17 170.22 ;
        RECT 0.5 170.22 14.24 170.29 ;
        RECT 0.5 170.29 14.31 170.36 ;
        RECT 0.5 170.36 14.38 170.43 ;
        RECT 0.5 170.43 14.45 170.5 ;
        RECT 0.5 170.5 14.52 170.57 ;
        RECT 0.5 170.57 14.59 170.64 ;
        RECT 0.5 170.64 14.66 170.71 ;
        RECT 0.5 170.71 14.73 170.78 ;
        RECT 0.5 170.78 14.8 170.85 ;
        RECT 0.5 170.85 14.87 170.92 ;
        RECT 0.5 170.92 14.94 170.99 ;
        RECT 0.5 164.68 13.96 169.94 ;
        RECT 0.5 163.63 14.94 163.7 ;
        RECT 0.5 163.7 14.87 163.77 ;
        RECT 0.5 163.77 14.8 163.84 ;
        RECT 0.5 163.84 14.73 163.91 ;
        RECT 0.5 163.91 14.66 163.98 ;
        RECT 0.5 163.98 14.59 164.05 ;
        RECT 0.5 164.05 14.52 164.12 ;
        RECT 0.5 164.12 14.45 164.19 ;
        RECT 0.5 164.19 14.38 164.26 ;
        RECT 0.5 164.26 14.31 164.33 ;
        RECT 0.5 164.33 14.24 164.4 ;
        RECT 0.5 164.4 14.17 164.47 ;
        RECT 0.5 164.47 14.1 164.54 ;
        RECT 0.5 164.54 14.03 164.61 ;
        RECT 0.5 164.61 13.96 164.68 ;
        RECT 0.5 160.99 68.01 163.63 ;
        RECT 0.5 159.94 13.96 160.01 ;
        RECT 0.5 160.01 14.03 160.08 ;
        RECT 0.5 160.08 14.1 160.15 ;
        RECT 0.5 160.15 14.17 160.22 ;
        RECT 0.5 160.22 14.24 160.29 ;
        RECT 0.5 160.29 14.31 160.36 ;
        RECT 0.5 160.36 14.38 160.43 ;
        RECT 0.5 160.43 14.45 160.5 ;
        RECT 0.5 160.5 14.52 160.57 ;
        RECT 0.5 160.57 14.59 160.64 ;
        RECT 0.5 160.64 14.66 160.71 ;
        RECT 0.5 160.71 14.73 160.78 ;
        RECT 0.5 160.78 14.8 160.85 ;
        RECT 0.5 160.85 14.87 160.92 ;
        RECT 0.5 160.92 14.94 160.99 ;
        RECT 0.5 154.68 13.96 159.94 ;
        RECT 0.5 153.63 14.94 153.7 ;
        RECT 0.5 153.7 14.87 153.77 ;
        RECT 0.5 153.77 14.8 153.84 ;
        RECT 0.5 153.84 14.73 153.91 ;
        RECT 0.5 153.91 14.66 153.98 ;
        RECT 0.5 153.98 14.59 154.05 ;
        RECT 0.5 154.05 14.52 154.12 ;
        RECT 0.5 154.12 14.45 154.19 ;
        RECT 0.5 154.19 14.38 154.26 ;
        RECT 0.5 154.26 14.31 154.33 ;
        RECT 0.5 154.33 14.24 154.4 ;
        RECT 0.5 154.4 14.17 154.47 ;
        RECT 0.5 154.47 14.1 154.54 ;
        RECT 0.5 154.54 14.03 154.61 ;
        RECT 0.5 154.61 13.96 154.68 ;
        RECT 0.5 150.99 68.01 153.63 ;
        RECT 0.5 149.94 13.96 150.01 ;
        RECT 0.5 150.01 14.03 150.08 ;
        RECT 0.5 150.08 14.1 150.15 ;
        RECT 0.5 150.15 14.17 150.22 ;
        RECT 0.5 150.22 14.24 150.29 ;
        RECT 0.5 150.29 14.31 150.36 ;
        RECT 0.5 150.36 14.38 150.43 ;
        RECT 0.5 150.43 14.45 150.5 ;
        RECT 0.5 150.5 14.52 150.57 ;
        RECT 0.5 150.57 14.59 150.64 ;
        RECT 0.5 150.64 14.66 150.71 ;
        RECT 0.5 150.71 14.73 150.78 ;
        RECT 0.5 150.78 14.8 150.85 ;
        RECT 0.5 150.85 14.87 150.92 ;
        RECT 0.5 150.92 14.94 150.99 ;
        RECT 0.5 144.68 13.96 149.94 ;
        RECT 0.5 143.63 14.94 143.7 ;
        RECT 0.5 143.7 14.87 143.77 ;
        RECT 0.5 143.77 14.8 143.84 ;
        RECT 0.5 143.84 14.73 143.91 ;
        RECT 0.5 143.91 14.66 143.98 ;
        RECT 0.5 143.98 14.59 144.05 ;
        RECT 0.5 144.05 14.52 144.12 ;
        RECT 0.5 144.12 14.45 144.19 ;
        RECT 0.5 144.19 14.38 144.26 ;
        RECT 0.5 144.26 14.31 144.33 ;
        RECT 0.5 144.33 14.24 144.4 ;
        RECT 0.5 144.4 14.17 144.47 ;
        RECT 0.5 144.47 14.1 144.54 ;
        RECT 0.5 144.54 14.03 144.61 ;
        RECT 0.5 144.61 13.96 144.68 ;
        RECT 0.5 140.99 68.01 143.63 ;
        RECT 0.5 139.94 13.96 140.01 ;
        RECT 0.5 140.01 14.03 140.08 ;
        RECT 0.5 140.08 14.1 140.15 ;
        RECT 0.5 140.15 14.17 140.22 ;
        RECT 0.5 140.22 14.24 140.29 ;
        RECT 0.5 140.29 14.31 140.36 ;
        RECT 0.5 140.36 14.38 140.43 ;
        RECT 0.5 140.43 14.45 140.5 ;
        RECT 0.5 140.5 14.52 140.57 ;
        RECT 0.5 140.57 14.59 140.64 ;
        RECT 0.5 140.64 14.66 140.71 ;
        RECT 0.5 140.71 14.73 140.78 ;
        RECT 0.5 140.78 14.8 140.85 ;
        RECT 0.5 140.85 14.87 140.92 ;
        RECT 0.5 140.92 14.94 140.99 ;
        RECT 0.5 134.68 13.96 139.94 ;
        RECT 0.5 133.63 14.94 133.7 ;
        RECT 0.5 133.7 14.87 133.77 ;
        RECT 0.5 133.77 14.8 133.84 ;
        RECT 0.5 133.84 14.73 133.91 ;
        RECT 0.5 133.91 14.66 133.98 ;
        RECT 0.5 133.98 14.59 134.05 ;
        RECT 0.5 134.05 14.52 134.12 ;
        RECT 0.5 134.12 14.45 134.19 ;
        RECT 0.5 134.19 14.38 134.26 ;
        RECT 0.5 134.26 14.31 134.33 ;
        RECT 0.5 134.33 14.24 134.4 ;
        RECT 0.5 134.4 14.17 134.47 ;
        RECT 0.5 134.47 14.1 134.54 ;
        RECT 0.5 134.54 14.03 134.61 ;
        RECT 0.5 134.61 13.96 134.68 ;
        RECT 0.5 130.99 68.01 133.63 ;
        RECT 0.5 129.94 13.96 130.01 ;
        RECT 0.5 130.01 14.03 130.08 ;
        RECT 0.5 130.08 14.1 130.15 ;
        RECT 0.5 130.15 14.17 130.22 ;
        RECT 0.5 130.22 14.24 130.29 ;
        RECT 0.5 130.29 14.31 130.36 ;
        RECT 0.5 130.36 14.38 130.43 ;
        RECT 0.5 130.43 14.45 130.5 ;
        RECT 0.5 130.5 14.52 130.57 ;
        RECT 0.5 130.57 14.59 130.64 ;
        RECT 0.5 130.64 14.66 130.71 ;
        RECT 0.5 130.71 14.73 130.78 ;
        RECT 0.5 130.78 14.8 130.85 ;
        RECT 0.5 130.85 14.87 130.92 ;
        RECT 0.5 130.92 14.94 130.99 ;
        RECT 0.5 124.68 13.96 129.94 ;
        RECT 0.5 123.14 15.43 123.21 ;
        RECT 0.5 123.21 15.36 123.28 ;
        RECT 0.5 123.28 15.29 123.35 ;
        RECT 0.5 123.35 15.22 123.42 ;
        RECT 0.5 123.42 15.15 123.49 ;
        RECT 0.5 123.49 15.08 123.56 ;
        RECT 0.5 123.56 15.01 123.63 ;
        RECT 0.5 123.63 14.94 123.7 ;
        RECT 0.5 123.7 14.87 123.77 ;
        RECT 0.5 123.77 14.8 123.84 ;
        RECT 0.5 123.84 14.73 123.91 ;
        RECT 0.5 123.91 14.66 123.98 ;
        RECT 0.5 123.98 14.59 124.05 ;
        RECT 0.5 124.05 14.52 124.12 ;
        RECT 0.5 124.12 14.45 124.19 ;
        RECT 0.5 124.19 14.38 124.26 ;
        RECT 0.5 124.26 14.31 124.33 ;
        RECT 0.5 124.33 14.24 124.4 ;
        RECT 0.5 124.4 14.17 124.47 ;
        RECT 0.5 124.47 14.1 124.54 ;
        RECT 0.5 124.54 14.03 124.61 ;
        RECT 0.5 124.61 13.96 124.68 ;
        RECT 0.5 76.045 15.5 123.14 ;
        RECT 0.5 74.295 13.75 74.365 ;
        RECT 0.5 74.365 13.82 74.435 ;
        RECT 0.5 74.435 13.89 74.505 ;
        RECT 0.5 74.505 13.96 74.575 ;
        RECT 0.5 74.575 14.03 74.645 ;
        RECT 0.5 74.645 14.1 74.715 ;
        RECT 0.5 74.715 14.17 74.785 ;
        RECT 0.5 74.785 14.24 74.855 ;
        RECT 0.5 74.855 14.31 74.925 ;
        RECT 0.5 74.925 14.38 74.995 ;
        RECT 0.5 74.995 14.45 75.065 ;
        RECT 0.5 75.065 14.52 75.135 ;
        RECT 0.5 75.135 14.59 75.205 ;
        RECT 0.5 75.205 14.66 75.275 ;
        RECT 0.5 75.275 14.73 75.345 ;
        RECT 0.5 75.345 14.8 75.415 ;
        RECT 0.5 75.415 14.87 75.485 ;
        RECT 0.5 75.485 14.94 75.555 ;
        RECT 0.5 75.555 15.01 75.625 ;
        RECT 0.5 75.625 15.08 75.695 ;
        RECT 0.5 75.695 15.15 75.765 ;
        RECT 0.5 75.765 15.22 75.835 ;
        RECT 0.5 75.835 15.29 75.905 ;
        RECT 0.5 75.905 15.36 75.975 ;
        RECT 0.5 75.975 15.43 76.045 ;
        RECT 0.5 24.165 13.75 74.295 ;
        RECT 0.5 24.16 13.75 24.165 ;
        RECT 0.5 24.09 13.755 24.16 ;
        RECT 0.5 24.02 13.825 24.09 ;
        RECT 0.5 23.95 13.895 24.02 ;
        RECT 0.5 23.88 13.965 23.95 ;
        RECT 0.5 23.81 14.035 23.88 ;
        RECT 0.5 23.74 14.105 23.81 ;
        RECT 0.5 23.67 14.175 23.74 ;
        RECT 0.5 23.6 14.245 23.67 ;
        RECT 0.5 23.53 14.315 23.6 ;
        RECT 0.5 23.46 14.385 23.53 ;
        RECT 0.5 23.39 14.455 23.46 ;
        RECT 0.5 23.32 14.525 23.39 ;
        RECT 0.5 23.25 14.595 23.32 ;
        RECT 0.5 23.18 14.665 23.25 ;
        RECT 0.5 23.11 14.735 23.18 ;
        RECT 0.5 23.04 14.805 23.11 ;
        RECT 0.5 22.97 14.875 23.04 ;
        RECT 0.5 22.9 14.945 22.97 ;
        RECT 0.5 22.83 15.015 22.9 ;
        RECT 0.5 22.76 15.085 22.83 ;
        RECT 0.5 22.69 15.155 22.76 ;
        RECT 0.5 22.62 15.225 22.69 ;
        RECT 0.5 22.55 15.295 22.62 ;
        RECT 0.5 22.48 15.365 22.55 ;
        RECT 0.5 22.41 15.435 22.48 ;
        RECT 0.5 22.34 15.505 22.41 ;
        RECT 0.5 22.27 15.575 22.34 ;
        RECT 0.5 22.2 15.645 22.27 ;
        RECT 0.5 22.13 15.715 22.2 ;
        RECT 0.5 22.06 15.785 22.13 ;
        RECT 0.5 21.99 15.855 22.06 ;
        RECT 0.5 21.92 15.925 21.99 ;
        RECT 0.5 21.85 15.995 21.92 ;
        RECT 0.5 21.78 16.065 21.85 ;
        RECT 0.5 21.71 16.135 21.78 ;
        RECT 0.5 21.64 16.205 21.71 ;
        RECT 0.5 21.57 16.275 21.64 ;
        RECT 0.5 21.5 16.345 21.57 ;
        RECT 0.5 21.43 16.415 21.5 ;
        RECT 0.5 21.36 16.485 21.43 ;
        RECT 0.5 21.29 16.555 21.36 ;
        RECT 0.5 21.22 16.625 21.29 ;
        RECT 0.5 21.15 16.695 21.22 ;
        RECT 0.5 21.08 16.765 21.15 ;
        RECT 0.5 21.01 16.835 21.08 ;
        RECT 0.5 20.94 16.905 21.01 ;
        RECT 0.5 20.87 16.975 20.94 ;
        RECT 0.5 20.8 17.045 20.87 ;
        RECT 0.5 20.73 17.115 20.8 ;
        RECT 0.5 20.66 17.185 20.73 ;
        RECT 0.5 20.59 17.255 20.66 ;
        RECT 0.5 20.52 17.325 20.59 ;
        RECT 0.5 20.45 17.395 20.52 ;
        RECT 0.5 20.38 17.465 20.45 ;
        RECT 0.5 20.31 17.535 20.38 ;
        RECT 0.5 20.24 17.605 20.31 ;
        RECT 0.5 20.17 17.675 20.24 ;
        RECT 0.5 20.1 17.745 20.17 ;
        RECT 0.5 20.03 17.815 20.1 ;
        RECT 0.5 19.96 17.885 20.03 ;
        RECT 0.5 19.89 17.955 19.96 ;
        RECT 0.5 19.82 18.025 19.89 ;
        RECT 0.5 19.75 18.095 19.82 ;
        RECT 0.5 19.68 18.165 19.75 ;
        RECT 0.5 19.61 18.235 19.68 ;
        RECT 0.5 19.54 18.305 19.61 ;
        RECT 0.5 19.47 18.375 19.54 ;
        RECT 0.5 19.4 18.445 19.47 ;
        RECT 0.5 19.33 18.515 19.4 ;
        RECT 0.5 19.26 18.585 19.33 ;
        RECT 0.5 19.19 18.655 19.26 ;
        RECT 0.5 19.12 18.725 19.19 ;
        RECT 0.5 19.05 18.795 19.12 ;
        RECT 0.5 18.98 18.865 19.05 ;
        RECT 0.5 18.91 18.935 18.98 ;
        RECT 0.5 18.84 19.005 18.91 ;
        RECT 0.5 18.77 19.075 18.84 ;
        RECT 0.5 18.7 19.145 18.77 ;
        RECT 0.5 18.63 19.215 18.7 ;
        RECT 0.5 18.56 19.285 18.63 ;
        RECT 0.5 18.49 19.355 18.56 ;
        RECT 0.5 18.42 19.425 18.49 ;
        RECT 0.5 18.35 19.495 18.42 ;
        RECT 0.5 18.28 19.565 18.35 ;
        RECT 0.5 18.21 19.635 18.28 ;
        RECT 0.5 18.14 19.705 18.21 ;
        RECT 0.5 18.07 19.775 18.14 ;
        RECT 0.5 18 19.845 18.07 ;
        RECT 0.5 17.93 19.915 18 ;
        RECT 0.5 17.86 19.985 17.93 ;
        RECT 0.5 17.79 20.055 17.86 ;
        RECT 0.5 17.72 20.125 17.79 ;
        RECT 0.5 17.65 20.195 17.72 ;
        RECT 0.5 17.58 20.265 17.65 ;
        RECT 0.5 17.51 20.335 17.58 ;
        RECT 0.5 17.44 20.405 17.51 ;
        RECT 0.5 17.37 20.475 17.44 ;
        RECT 0.5 17.3 20.545 17.37 ;
        RECT 0.5 17.23 20.615 17.3 ;
        RECT 0.5 17.16 20.685 17.23 ;
        RECT 0.5 17.09 20.755 17.16 ;
        RECT 0.5 17.02 20.825 17.09 ;
        RECT 0.5 16.95 20.895 17.02 ;
        RECT 0.5 16.88 20.965 16.95 ;
        RECT 0.5 16.81 21.035 16.88 ;
        RECT 0.5 16.74 21.105 16.81 ;
        RECT 0.5 16.67 21.175 16.74 ;
        RECT 0.5 16.6 21.245 16.67 ;
        RECT 0.5 16.53 21.315 16.6 ;
        RECT 0.5 16.46 21.385 16.53 ;
        RECT 0.5 16.39 21.455 16.46 ;
        RECT 0.5 16.32 21.525 16.39 ;
        RECT 0.5 16.25 21.595 16.32 ;
        RECT 0.5 16.18 21.665 16.25 ;
        RECT 0.5 9.18 55.595 16.18 ;
        RECT 0.5 9.105 17.5 9.14 ;
        RECT 0.5 9.14 17.535 9.175 ;
        RECT 0.5 9.175 17.57 9.18 ;
        RECT 12.015 8.72 17.115 8.79 ;
        RECT 11.945 8.79 17.185 8.86 ;
        RECT 11.875 8.86 17.255 8.93 ;
        RECT 11.805 8.93 17.325 9 ;
        RECT 11.735 9 17.395 9.07 ;
        RECT 11.665 9.07 17.465 9.105 ;
        RECT 0.5 8.71 10.42 8.78 ;
        RECT 0.5 8.78 10.49 8.85 ;
        RECT 0.5 8.85 10.56 8.92 ;
        RECT 0.5 8.92 10.63 8.99 ;
        RECT 0.5 8.99 10.7 9.06 ;
        RECT 0.5 9.06 10.77 9.105 ;
        RECT 12.015 8.465 16.86 8.535 ;
        RECT 12.015 8.535 16.93 8.605 ;
        RECT 12.015 8.605 17 8.675 ;
        RECT 12.015 8.675 17.07 8.72 ;
        RECT 0.5 6.94 10.42 8.71 ;
        RECT 12.015 6.935 16.86 8.465 ;
        RECT 0.5 6.545 10.745 6.615 ;
        RECT 0.5 6.615 10.675 6.685 ;
        RECT 0.5 6.685 10.605 6.755 ;
        RECT 0.5 6.755 10.535 6.825 ;
        RECT 0.5 6.825 10.465 6.895 ;
        RECT 0.5 6.895 10.42 6.94 ;
        RECT 11.695 6.545 16.86 6.615 ;
        RECT 11.765 6.615 16.86 6.685 ;
        RECT 11.835 6.685 16.86 6.755 ;
        RECT 11.905 6.755 16.86 6.825 ;
        RECT 11.975 6.825 16.86 6.895 ;
        RECT 12.015 6.895 16.86 6.935 ;
        RECT 0.5 4.21 16.86 6.545 ;
        RECT 0.5 0.575 20.425 0.645 ;
        RECT 0.5 0.645 20.355 0.715 ;
        RECT 0.5 0.715 20.285 0.785 ;
        RECT 0.5 0.785 20.215 0.855 ;
        RECT 0.5 0.855 20.145 0.925 ;
        RECT 0.5 0.925 20.075 0.995 ;
        RECT 0.5 0.995 20.005 1.065 ;
        RECT 0.5 1.065 19.935 1.135 ;
        RECT 0.5 1.135 19.865 1.205 ;
        RECT 0.5 1.205 19.795 1.275 ;
        RECT 0.5 1.275 19.725 1.345 ;
        RECT 0.5 1.345 19.655 1.415 ;
        RECT 0.5 1.415 19.585 1.485 ;
        RECT 0.5 1.485 19.515 1.555 ;
        RECT 0.5 1.555 19.445 1.625 ;
        RECT 0.5 1.625 19.375 1.695 ;
        RECT 0.5 1.695 19.305 1.765 ;
        RECT 0.5 1.765 19.235 1.835 ;
        RECT 0.5 1.835 19.165 1.905 ;
        RECT 0.5 1.905 19.095 1.975 ;
        RECT 0.5 1.975 19.025 2.045 ;
        RECT 0.5 2.045 18.955 2.115 ;
        RECT 0.5 2.115 18.885 2.185 ;
        RECT 0.5 2.185 18.815 2.255 ;
        RECT 0.5 2.255 18.745 2.325 ;
        RECT 0.5 2.325 18.675 2.395 ;
        RECT 0.5 2.395 18.605 2.465 ;
        RECT 0.5 2.465 18.535 2.535 ;
        RECT 0.5 2.535 18.465 2.605 ;
        RECT 0.5 2.605 18.395 2.675 ;
        RECT 0.5 2.675 18.325 2.745 ;
        RECT 0.5 2.745 18.255 2.815 ;
        RECT 0.5 2.815 18.185 2.885 ;
        RECT 0.5 2.885 18.115 2.955 ;
        RECT 0.5 2.955 18.045 3.025 ;
        RECT 0.5 3.025 17.975 3.095 ;
        RECT 0.5 3.095 17.905 3.165 ;
        RECT 0.5 3.165 17.835 3.235 ;
        RECT 0.5 3.235 17.765 3.305 ;
        RECT 0.5 3.305 17.695 3.375 ;
        RECT 0.5 3.375 17.625 3.445 ;
        RECT 0.5 3.445 17.555 3.515 ;
        RECT 0.5 3.515 17.485 3.585 ;
        RECT 0.5 3.585 17.415 3.655 ;
        RECT 0.5 3.655 17.345 3.725 ;
        RECT 0.5 3.725 17.275 3.795 ;
        RECT 0.5 3.795 17.205 3.865 ;
        RECT 0.5 3.865 17.135 3.935 ;
        RECT 0.5 3.935 17.065 4.005 ;
        RECT 0.5 4.005 16.995 4.075 ;
        RECT 0.5 4.075 16.925 4.145 ;
        RECT 0.5 4.145 16.86 4.21 ;
        RECT 0.5 0 20.495 0.575 ;
    END
  END src_bdy_lvc1

  PIN ogc_lvc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 25.04 0 25.46 24.385 ;
    END
  END ogc_lvc

  PIN drn_lvc1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605 170.61 25.115 189.515 ;
        RECT 37.945 169.025 48.835 189.515 ;
        RECT 49.87 168.92 60.33 189.515 ;
        RECT 26.035 167.46 36.925 189.515 ;
        RECT 15.605 167.1 21.605 167.25 ;
        RECT 15.605 167.25 21.755 167.4 ;
        RECT 15.605 167.4 21.905 167.55 ;
        RECT 15.605 167.55 22.055 167.7 ;
        RECT 15.605 167.7 22.205 167.85 ;
        RECT 15.605 167.85 22.355 168 ;
        RECT 15.605 168 22.505 168.15 ;
        RECT 15.605 168.15 22.655 168.3 ;
        RECT 15.605 168.3 22.805 168.45 ;
        RECT 15.605 168.45 22.955 168.6 ;
        RECT 15.605 168.6 23.105 168.75 ;
        RECT 15.605 168.75 23.255 168.9 ;
        RECT 15.605 168.9 23.405 169.05 ;
        RECT 15.605 169.05 23.555 169.2 ;
        RECT 15.605 169.2 23.705 169.35 ;
        RECT 15.605 169.35 23.855 169.5 ;
        RECT 15.605 169.5 24.005 169.65 ;
        RECT 15.605 169.65 24.155 169.8 ;
        RECT 15.605 169.8 24.305 169.95 ;
        RECT 15.605 169.95 24.455 170.1 ;
        RECT 15.605 170.1 24.605 170.25 ;
        RECT 15.605 170.25 24.755 170.4 ;
        RECT 15.605 170.4 24.905 170.55 ;
        RECT 15.605 170.55 25.055 170.61 ;
        RECT 54.33 164.46 60.33 164.61 ;
        RECT 54.18 164.61 60.33 164.76 ;
        RECT 54.03 164.76 60.33 164.91 ;
        RECT 53.88 164.91 60.33 165.06 ;
        RECT 53.73 165.06 60.33 165.21 ;
        RECT 53.58 165.21 60.33 165.36 ;
        RECT 53.43 165.36 60.33 165.51 ;
        RECT 53.28 165.51 60.33 165.66 ;
        RECT 53.13 165.66 60.33 165.81 ;
        RECT 52.98 165.81 60.33 165.96 ;
        RECT 52.83 165.96 60.33 166.11 ;
        RECT 52.68 166.11 60.33 166.26 ;
        RECT 52.53 166.26 60.33 166.41 ;
        RECT 52.38 166.41 60.33 166.56 ;
        RECT 52.23 166.56 60.33 166.71 ;
        RECT 52.08 166.71 60.33 166.86 ;
        RECT 51.93 166.86 60.33 167.01 ;
        RECT 51.78 167.01 60.33 167.16 ;
        RECT 51.63 167.16 60.33 167.31 ;
        RECT 51.48 167.31 60.33 167.46 ;
        RECT 51.33 167.46 60.33 167.61 ;
        RECT 51.18 167.61 60.33 167.76 ;
        RECT 51.03 167.76 60.33 167.91 ;
        RECT 50.88 167.91 60.33 168.06 ;
        RECT 50.73 168.06 60.33 168.21 ;
        RECT 50.58 168.21 60.33 168.36 ;
        RECT 50.43 168.36 60.33 168.51 ;
        RECT 50.28 168.51 60.33 168.66 ;
        RECT 50.13 168.66 60.33 168.81 ;
        RECT 49.98 168.81 60.33 168.92 ;
        RECT 42.835 164.135 48.835 164.285 ;
        RECT 42.685 164.285 48.835 164.435 ;
        RECT 42.535 164.435 48.835 164.585 ;
        RECT 42.385 164.585 48.835 164.735 ;
        RECT 42.235 164.735 48.835 164.885 ;
        RECT 42.085 164.885 48.835 165.035 ;
        RECT 41.935 165.035 48.835 165.185 ;
        RECT 41.785 165.185 48.835 165.335 ;
        RECT 41.635 165.335 48.835 165.485 ;
        RECT 41.485 165.485 48.835 165.635 ;
        RECT 41.335 165.635 48.835 165.785 ;
        RECT 41.185 165.785 48.835 165.935 ;
        RECT 41.035 165.935 48.835 166.085 ;
        RECT 40.885 166.085 48.835 166.235 ;
        RECT 40.735 166.235 48.835 166.385 ;
        RECT 40.585 166.385 48.835 166.535 ;
        RECT 40.435 166.535 48.835 166.685 ;
        RECT 40.285 166.685 48.835 166.835 ;
        RECT 40.135 166.835 48.835 166.985 ;
        RECT 39.985 166.985 48.835 167.135 ;
        RECT 39.835 167.135 48.835 167.285 ;
        RECT 39.685 167.285 48.835 167.435 ;
        RECT 39.535 167.435 48.835 167.585 ;
        RECT 39.385 167.585 48.835 167.735 ;
        RECT 39.235 167.735 48.835 167.885 ;
        RECT 39.085 167.885 48.835 168.035 ;
        RECT 38.935 168.035 48.835 168.185 ;
        RECT 38.785 168.185 48.835 168.335 ;
        RECT 38.635 168.335 48.835 168.485 ;
        RECT 38.485 168.485 48.835 168.635 ;
        RECT 38.335 168.635 48.835 168.785 ;
        RECT 38.185 168.785 48.835 168.935 ;
        RECT 38.035 168.935 48.835 169.025 ;
        RECT 26.035 162.57 32.035 162.72 ;
        RECT 26.035 162.72 32.185 162.87 ;
        RECT 26.035 162.87 32.335 163.02 ;
        RECT 26.035 163.02 32.485 163.17 ;
        RECT 26.035 163.17 32.635 163.32 ;
        RECT 26.035 163.32 32.785 163.47 ;
        RECT 26.035 163.47 32.935 163.62 ;
        RECT 26.035 163.62 33.085 163.77 ;
        RECT 26.035 163.77 33.235 163.92 ;
        RECT 26.035 163.92 33.385 164.07 ;
        RECT 26.035 164.07 33.535 164.22 ;
        RECT 26.035 164.22 33.685 164.37 ;
        RECT 26.035 164.37 33.835 164.52 ;
        RECT 26.035 164.52 33.985 164.67 ;
        RECT 26.035 164.67 34.135 164.82 ;
        RECT 26.035 164.82 34.285 164.97 ;
        RECT 26.035 164.97 34.435 165.12 ;
        RECT 26.035 165.12 34.585 165.27 ;
        RECT 26.035 165.27 34.735 165.42 ;
        RECT 26.035 165.42 34.885 165.57 ;
        RECT 26.035 165.57 35.035 165.72 ;
        RECT 26.035 165.72 35.185 165.87 ;
        RECT 26.035 165.87 35.335 166.02 ;
        RECT 26.035 166.02 35.485 166.17 ;
        RECT 26.035 166.17 35.635 166.32 ;
        RECT 26.035 166.32 35.785 166.47 ;
        RECT 26.035 166.47 35.935 166.62 ;
        RECT 26.035 166.62 36.085 166.77 ;
        RECT 26.035 166.77 36.235 166.92 ;
        RECT 26.035 166.92 36.385 167.07 ;
        RECT 26.035 167.07 36.535 167.22 ;
        RECT 26.035 167.22 36.685 167.37 ;
        RECT 26.035 167.37 36.835 167.46 ;
        RECT 54.33 100.165 60.33 164.46 ;
        RECT 52 97.685 60.33 97.835 ;
        RECT 52.15 97.835 60.33 97.985 ;
        RECT 52.3 97.985 60.33 98.135 ;
        RECT 52.45 98.135 60.33 98.285 ;
        RECT 52.6 98.285 60.33 98.435 ;
        RECT 52.75 98.435 60.33 98.585 ;
        RECT 52.9 98.585 60.33 98.735 ;
        RECT 53.05 98.735 60.33 98.885 ;
        RECT 53.2 98.885 60.33 99.035 ;
        RECT 53.35 99.035 60.33 99.185 ;
        RECT 53.5 99.185 60.33 99.335 ;
        RECT 53.65 99.335 60.33 99.485 ;
        RECT 53.8 99.485 60.33 99.635 ;
        RECT 53.95 99.635 60.33 99.785 ;
        RECT 54.1 99.785 60.33 99.935 ;
        RECT 54.25 99.935 60.33 100.085 ;
        RECT 54.33 100.085 60.33 100.165 ;
        RECT 42.835 96.81 48.835 164.135 ;
        RECT 15.605 96.79 21.605 167.1 ;
        RECT 42.835 95.415 47.44 95.565 ;
        RECT 42.835 95.565 47.59 95.715 ;
        RECT 42.835 95.715 47.74 95.865 ;
        RECT 42.835 95.865 47.89 96.015 ;
        RECT 42.835 96.015 48.04 96.165 ;
        RECT 42.835 96.165 48.19 96.315 ;
        RECT 42.835 96.315 48.34 96.465 ;
        RECT 42.835 96.465 48.49 96.615 ;
        RECT 42.835 96.615 48.64 96.765 ;
        RECT 42.835 96.765 48.79 96.81 ;
        RECT 26.035 94.5 32.035 162.57 ;
        RECT 15.605 94.31 23.935 94.46 ;
        RECT 15.605 94.46 23.785 94.61 ;
        RECT 15.605 94.61 23.635 94.76 ;
        RECT 15.605 94.76 23.485 94.91 ;
        RECT 15.605 94.91 23.335 95.06 ;
        RECT 15.605 95.06 23.185 95.21 ;
        RECT 15.605 95.21 23.035 95.36 ;
        RECT 15.605 95.36 22.885 95.51 ;
        RECT 15.605 95.51 22.735 95.66 ;
        RECT 15.605 95.66 22.585 95.81 ;
        RECT 15.605 95.81 22.435 95.96 ;
        RECT 15.605 95.96 22.285 96.11 ;
        RECT 15.605 96.11 22.135 96.26 ;
        RECT 15.605 96.26 21.985 96.41 ;
        RECT 15.605 96.41 21.835 96.56 ;
        RECT 15.605 96.56 21.685 96.71 ;
        RECT 15.605 96.71 21.605 96.79 ;
        RECT 27.145 93.39 32.035 93.54 ;
        RECT 26.995 93.54 32.035 93.69 ;
        RECT 26.845 93.69 32.035 93.84 ;
        RECT 26.695 93.84 32.035 93.99 ;
        RECT 26.545 93.99 32.035 94.14 ;
        RECT 26.395 94.14 32.035 94.29 ;
        RECT 26.245 94.29 32.035 94.44 ;
        RECT 26.095 94.44 32.035 94.5 ;
        RECT 37.945 90.375 42.4 90.525 ;
        RECT 38.095 90.525 42.55 90.675 ;
        RECT 38.245 90.675 42.7 90.825 ;
        RECT 38.395 90.825 42.85 90.975 ;
        RECT 38.545 90.975 43 91.125 ;
        RECT 38.695 91.125 43.15 91.275 ;
        RECT 38.845 91.275 43.3 91.425 ;
        RECT 38.995 91.425 43.45 91.575 ;
        RECT 39.145 91.575 43.6 91.725 ;
        RECT 39.295 91.725 43.75 91.875 ;
        RECT 39.445 91.875 43.9 92.025 ;
        RECT 39.595 92.025 44.05 92.175 ;
        RECT 39.745 92.175 44.2 92.325 ;
        RECT 39.895 92.325 44.35 92.475 ;
        RECT 40.045 92.475 44.5 92.625 ;
        RECT 40.195 92.625 44.65 92.775 ;
        RECT 40.345 92.775 44.8 92.925 ;
        RECT 40.495 92.925 44.95 93.075 ;
        RECT 40.645 93.075 45.1 93.225 ;
        RECT 40.795 93.225 45.25 93.375 ;
        RECT 40.945 93.375 45.4 93.525 ;
        RECT 41.095 93.525 45.55 93.675 ;
        RECT 41.245 93.675 45.7 93.825 ;
        RECT 41.395 93.825 45.85 93.975 ;
        RECT 41.545 93.975 46 94.125 ;
        RECT 41.695 94.125 46.15 94.275 ;
        RECT 41.845 94.275 46.3 94.425 ;
        RECT 41.995 94.425 46.45 94.575 ;
        RECT 42.145 94.575 46.6 94.725 ;
        RECT 42.295 94.725 46.75 94.875 ;
        RECT 42.445 94.875 46.9 95.025 ;
        RECT 42.595 95.025 47.05 95.175 ;
        RECT 42.745 95.175 47.2 95.325 ;
        RECT 42.835 95.325 47.35 95.415 ;
        RECT 30.16 90.375 34.9 90.525 ;
        RECT 30.01 90.525 34.75 90.675 ;
        RECT 29.86 90.675 34.6 90.825 ;
        RECT 29.71 90.825 34.45 90.975 ;
        RECT 29.56 90.975 34.3 91.125 ;
        RECT 29.41 91.125 34.15 91.275 ;
        RECT 29.26 91.275 34 91.425 ;
        RECT 29.11 91.425 33.85 91.575 ;
        RECT 28.96 91.575 33.7 91.725 ;
        RECT 28.81 91.725 33.55 91.875 ;
        RECT 28.66 91.875 33.4 92.025 ;
        RECT 28.51 92.025 33.25 92.175 ;
        RECT 28.36 92.175 33.1 92.325 ;
        RECT 28.21 92.325 32.95 92.475 ;
        RECT 28.06 92.475 32.8 92.625 ;
        RECT 27.91 92.625 32.65 92.775 ;
        RECT 27.76 92.775 32.5 92.925 ;
        RECT 27.61 92.925 32.35 93.075 ;
        RECT 27.46 93.075 32.2 93.225 ;
        RECT 27.31 93.225 32.05 93.375 ;
        RECT 27.16 93.375 32.035 93.39 ;
        RECT 42.69 88.375 51.02 88.525 ;
        RECT 42.84 88.525 51.17 88.675 ;
        RECT 42.99 88.675 51.32 88.825 ;
        RECT 43.14 88.825 51.47 88.975 ;
        RECT 43.29 88.975 51.62 89.125 ;
        RECT 43.44 89.125 51.77 89.275 ;
        RECT 43.59 89.275 51.92 89.425 ;
        RECT 43.74 89.425 52.07 89.575 ;
        RECT 43.89 89.575 52.22 89.725 ;
        RECT 44.04 89.725 52.37 89.875 ;
        RECT 44.19 89.875 52.52 90.025 ;
        RECT 44.34 90.025 52.67 90.175 ;
        RECT 44.49 90.175 52.82 90.325 ;
        RECT 44.64 90.325 52.97 90.475 ;
        RECT 44.79 90.475 53.12 90.625 ;
        RECT 44.94 90.625 53.27 90.775 ;
        RECT 45.09 90.775 53.42 90.925 ;
        RECT 45.24 90.925 53.57 91.075 ;
        RECT 45.39 91.075 53.72 91.225 ;
        RECT 45.54 91.225 53.87 91.375 ;
        RECT 45.69 91.375 54.02 91.525 ;
        RECT 45.84 91.525 54.17 91.675 ;
        RECT 45.99 91.675 54.32 91.825 ;
        RECT 46.14 91.825 54.47 91.975 ;
        RECT 46.29 91.975 54.62 92.125 ;
        RECT 46.44 92.125 54.77 92.275 ;
        RECT 46.59 92.275 54.92 92.425 ;
        RECT 46.74 92.425 55.07 92.575 ;
        RECT 46.89 92.575 55.22 92.725 ;
        RECT 47.04 92.725 55.37 92.875 ;
        RECT 47.19 92.875 55.52 93.025 ;
        RECT 47.34 93.025 55.67 93.175 ;
        RECT 47.49 93.175 55.82 93.325 ;
        RECT 47.64 93.325 55.97 93.475 ;
        RECT 47.79 93.475 56.12 93.625 ;
        RECT 47.94 93.625 56.27 93.775 ;
        RECT 48.09 93.775 56.42 93.925 ;
        RECT 48.24 93.925 56.57 94.075 ;
        RECT 48.39 94.075 56.72 94.225 ;
        RECT 48.54 94.225 56.87 94.375 ;
        RECT 48.69 94.375 57.02 94.525 ;
        RECT 48.84 94.525 57.17 94.675 ;
        RECT 48.99 94.675 57.32 94.825 ;
        RECT 49.14 94.825 57.47 94.975 ;
        RECT 49.29 94.975 57.62 95.125 ;
        RECT 49.44 95.125 57.77 95.275 ;
        RECT 49.59 95.275 57.92 95.425 ;
        RECT 49.74 95.425 58.07 95.575 ;
        RECT 49.89 95.575 58.22 95.725 ;
        RECT 50.04 95.725 58.37 95.875 ;
        RECT 50.19 95.875 58.52 96.025 ;
        RECT 50.34 96.025 58.67 96.175 ;
        RECT 50.49 96.175 58.82 96.325 ;
        RECT 50.64 96.325 58.97 96.475 ;
        RECT 50.79 96.475 59.12 96.625 ;
        RECT 50.94 96.625 59.27 96.775 ;
        RECT 51.09 96.775 59.42 96.925 ;
        RECT 51.24 96.925 59.57 97.075 ;
        RECT 51.39 97.075 59.72 97.225 ;
        RECT 51.54 97.225 59.87 97.375 ;
        RECT 51.69 97.375 60.02 97.525 ;
        RECT 51.84 97.525 60.17 97.675 ;
        RECT 51.85 97.675 60.32 97.685 ;
        RECT 41.76 87.445 51.02 87.595 ;
        RECT 41.91 87.595 51.02 87.745 ;
        RECT 42.06 87.745 51.02 87.895 ;
        RECT 42.21 87.895 51.02 88.045 ;
        RECT 42.36 88.045 51.02 88.195 ;
        RECT 42.51 88.195 51.02 88.345 ;
        RECT 42.54 88.345 51.02 88.375 ;
        RECT 33.175 87.36 39.385 87.51 ;
        RECT 33.025 87.51 39.535 87.66 ;
        RECT 32.875 87.66 39.685 87.81 ;
        RECT 32.725 87.81 39.835 87.96 ;
        RECT 32.575 87.96 39.985 88.11 ;
        RECT 32.425 88.11 40.135 88.26 ;
        RECT 32.275 88.26 40.285 88.41 ;
        RECT 32.125 88.41 40.435 88.56 ;
        RECT 31.975 88.56 40.585 88.71 ;
        RECT 31.825 88.71 40.735 88.86 ;
        RECT 31.675 88.86 40.885 89.01 ;
        RECT 31.525 89.01 41.035 89.16 ;
        RECT 31.375 89.16 41.185 89.31 ;
        RECT 31.225 89.31 41.335 89.46 ;
        RECT 31.075 89.46 41.485 89.61 ;
        RECT 30.925 89.61 41.635 89.76 ;
        RECT 30.775 89.76 41.785 89.91 ;
        RECT 30.625 89.91 41.935 90.06 ;
        RECT 30.475 90.06 42.085 90.21 ;
        RECT 30.325 90.21 42.235 90.36 ;
        RECT 30.175 90.36 42.385 90.375 ;
        RECT 41.61 86.96 51.02 87.445 ;
        RECT 23.665 86.25 31.995 86.4 ;
        RECT 23.515 86.4 31.845 86.55 ;
        RECT 23.365 86.55 31.695 86.7 ;
        RECT 23.215 86.7 31.545 86.85 ;
        RECT 23.065 86.85 31.395 87 ;
        RECT 22.915 87 31.245 87.15 ;
        RECT 22.765 87.15 31.095 87.3 ;
        RECT 22.615 87.3 30.945 87.45 ;
        RECT 22.465 87.45 30.795 87.6 ;
        RECT 22.315 87.6 30.645 87.75 ;
        RECT 22.165 87.75 30.495 87.9 ;
        RECT 22.015 87.9 30.345 88.05 ;
        RECT 21.865 88.05 30.195 88.2 ;
        RECT 21.715 88.2 30.045 88.35 ;
        RECT 21.565 88.35 29.895 88.5 ;
        RECT 21.415 88.5 29.745 88.65 ;
        RECT 21.265 88.65 29.595 88.8 ;
        RECT 21.115 88.8 29.445 88.95 ;
        RECT 20.965 88.95 29.295 89.1 ;
        RECT 20.815 89.1 29.145 89.25 ;
        RECT 20.665 89.25 28.995 89.4 ;
        RECT 20.515 89.4 28.845 89.55 ;
        RECT 20.365 89.55 28.695 89.7 ;
        RECT 20.215 89.7 28.545 89.85 ;
        RECT 20.065 89.85 28.395 90 ;
        RECT 19.915 90 28.245 90.15 ;
        RECT 19.765 90.15 28.095 90.3 ;
        RECT 19.615 90.3 27.945 90.45 ;
        RECT 19.465 90.45 27.795 90.6 ;
        RECT 19.315 90.6 27.645 90.75 ;
        RECT 19.165 90.75 27.495 90.9 ;
        RECT 19.015 90.9 27.345 91.05 ;
        RECT 18.865 91.05 27.195 91.2 ;
        RECT 18.715 91.2 27.045 91.35 ;
        RECT 18.565 91.35 26.895 91.5 ;
        RECT 18.415 91.5 26.745 91.65 ;
        RECT 18.265 91.65 26.595 91.8 ;
        RECT 18.115 91.8 26.445 91.95 ;
        RECT 17.965 91.95 26.295 92.1 ;
        RECT 17.815 92.1 26.145 92.25 ;
        RECT 17.665 92.25 25.995 92.4 ;
        RECT 17.515 92.4 25.845 92.55 ;
        RECT 17.365 92.55 25.695 92.7 ;
        RECT 17.215 92.7 25.545 92.85 ;
        RECT 17.065 92.85 25.395 93 ;
        RECT 16.915 93 25.245 93.15 ;
        RECT 16.765 93.15 25.095 93.3 ;
        RECT 16.615 93.3 24.945 93.45 ;
        RECT 16.465 93.45 24.795 93.6 ;
        RECT 16.315 93.6 24.645 93.75 ;
        RECT 16.165 93.75 24.495 93.9 ;
        RECT 16.015 93.9 24.345 94.05 ;
        RECT 15.865 94.05 24.195 94.2 ;
        RECT 15.715 94.2 24.085 94.31 ;
        RECT 23.85 86.065 32.145 86.155 ;
        RECT 23.76 86.155 32.145 86.245 ;
        RECT 23.67 86.245 32.145 86.25 ;
        RECT 34.505 86.03 39.385 86.18 ;
        RECT 34.355 86.18 39.385 86.33 ;
        RECT 34.205 86.33 39.385 86.48 ;
        RECT 34.055 86.48 39.385 86.63 ;
        RECT 33.905 86.63 39.385 86.78 ;
        RECT 33.755 86.78 39.385 86.93 ;
        RECT 33.605 86.93 39.385 87.08 ;
        RECT 33.455 87.08 39.385 87.23 ;
        RECT 33.305 87.23 39.385 87.36 ;
        RECT 41.61 84.81 48.87 84.96 ;
        RECT 41.61 84.96 49.02 85.11 ;
        RECT 41.61 85.11 49.17 85.26 ;
        RECT 41.61 85.26 49.32 85.41 ;
        RECT 41.61 85.41 49.47 85.56 ;
        RECT 41.61 85.56 49.62 85.71 ;
        RECT 41.61 85.71 49.77 85.86 ;
        RECT 41.61 85.86 49.92 86.01 ;
        RECT 41.61 86.01 50.07 86.16 ;
        RECT 41.61 86.16 50.22 86.31 ;
        RECT 41.61 86.31 50.37 86.46 ;
        RECT 41.61 86.46 50.52 86.61 ;
        RECT 41.61 86.61 50.67 86.76 ;
        RECT 41.61 86.76 50.82 86.91 ;
        RECT 41.61 86.91 50.97 86.96 ;
        RECT 23.85 84.69 32.145 86.065 ;
        RECT 34.505 84.69 39.385 86.03 ;
        RECT 41.61 84.69 48.87 84.81 ;
        RECT 23.85 84.65 32.165 84.67 ;
        RECT 23.85 84.67 32.145 84.69 ;
        RECT 33.945 83.98 39.945 84.13 ;
        RECT 34.095 84.13 39.795 84.28 ;
        RECT 34.245 84.28 39.645 84.43 ;
        RECT 34.395 84.43 39.495 84.58 ;
        RECT 34.505 84.58 39.385 84.69 ;
        RECT 41.05 83.98 48.87 84.13 ;
        RECT 41.2 84.13 48.87 84.28 ;
        RECT 41.35 84.28 48.87 84.43 ;
        RECT 41.5 84.43 48.87 84.58 ;
        RECT 41.61 84.58 48.87 84.69 ;
        RECT 24.52 83.98 32.705 84.13 ;
        RECT 24.37 84.13 32.555 84.28 ;
        RECT 24.22 84.28 32.405 84.43 ;
        RECT 24.07 84.43 32.255 84.58 ;
        RECT 23.92 84.58 32.185 84.65 ;
        RECT 26 82.5 48.87 82.65 ;
        RECT 25.85 82.65 48.87 82.8 ;
        RECT 25.7 82.8 48.87 82.95 ;
        RECT 25.55 82.95 48.87 83.1 ;
        RECT 25.4 83.1 48.87 83.25 ;
        RECT 25.25 83.25 48.87 83.4 ;
        RECT 25.1 83.4 48.87 83.55 ;
        RECT 24.95 83.55 48.87 83.7 ;
        RECT 24.8 83.7 48.87 83.85 ;
        RECT 24.65 83.85 48.87 83.98 ;
        RECT 26 76.815 48.87 82.5 ;
        RECT 26 74.74 46.795 74.89 ;
        RECT 26 74.89 46.945 75.04 ;
        RECT 26 75.04 47.095 75.19 ;
        RECT 26 75.19 47.245 75.34 ;
        RECT 26 75.34 47.395 75.49 ;
        RECT 26 75.49 47.545 75.64 ;
        RECT 26 75.64 47.695 75.79 ;
        RECT 26 75.79 47.845 75.94 ;
        RECT 26 75.94 47.995 76.09 ;
        RECT 26 76.09 48.145 76.24 ;
        RECT 26 76.24 48.295 76.39 ;
        RECT 26 76.39 48.445 76.54 ;
        RECT 26 76.54 48.595 76.69 ;
        RECT 26 76.69 48.745 76.815 ;
        RECT 26 71.105 36.88 71.255 ;
        RECT 26 71.255 37.03 71.405 ;
        RECT 26 71.405 37.18 71.555 ;
        RECT 26 71.555 37.33 71.705 ;
        RECT 26 71.705 37.48 71.855 ;
        RECT 26 71.855 37.63 72.005 ;
        RECT 26 72.005 37.78 72.155 ;
        RECT 26 72.155 37.93 72.305 ;
        RECT 26 72.305 38.08 72.455 ;
        RECT 26 72.455 38.23 72.605 ;
        RECT 26 72.605 38.38 72.755 ;
        RECT 26 72.755 38.53 72.905 ;
        RECT 26 72.905 38.68 73.055 ;
        RECT 26 73.055 38.83 73.205 ;
        RECT 26 73.205 38.98 73.355 ;
        RECT 26 73.355 39.13 73.505 ;
        RECT 26 73.505 39.28 73.655 ;
        RECT 26 73.655 39.43 73.805 ;
        RECT 26 73.805 39.58 73.955 ;
        RECT 26 73.955 39.73 74.105 ;
        RECT 26 74.105 39.88 74.255 ;
        RECT 26 74.255 40.03 74.405 ;
        RECT 26 74.405 40.18 74.555 ;
        RECT 26 74.555 40.33 74.705 ;
        RECT 26 74.705 40.48 74.74 ;
        RECT 26 0 36.88 71.105 ;
    END
  END drn_lvc1

  PIN drn_lvc2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.38 0 49.255 69.49 ;
    END
  END drn_lvc2
  OBS
    LAYER met2 ;
      RECT 14.24 144.795 75 149.825 ;
      RECT 15.125 143.91 75 144.795 ;
      RECT 15.66 143.77 75 143.91 ;
      RECT 68.15 140.85 75 143.77 ;
      RECT 15.52 140.71 75 140.85 ;
      RECT 14.24 139.825 75 140.71 ;
      RECT 14.24 134.795 75 139.825 ;
      RECT 15.125 133.91 75 134.795 ;
      RECT 15.66 133.77 75 133.91 ;
      RECT 68.15 130.85 75 133.77 ;
      RECT 15.52 130.71 75 130.85 ;
      RECT 14.24 129.825 75 130.71 ;
      RECT 14.24 124.795 75 129.825 ;
      RECT 15.78 123.255 75 124.795 ;
      RECT 15.78 98.7 75 123.255 ;
      RECT 15.78 75.93 65.86 98.7 ;
      RECT 68.15 74.49 75 98.7 ;
      RECT 14.34 74.49 65.86 75.93 ;
      RECT 14.03 74.18 65.86 74.49 ;
      RECT 68.865 73.77 75 74.49 ;
      RECT 14.03 73.77 65.55 74.18 ;
      RECT 14.03 70.85 15.995 73.77 ;
      RECT 14.03 69.88 64.885 70.85 ;
      RECT 14.03 64.735 65.855 69.88 ;
      RECT 14.03 63.77 65.855 64.735 ;
      RECT 14.03 60.85 15.995 63.77 ;
      RECT 14.03 59.88 64.885 60.85 ;
      RECT 14.03 54.745 65.855 59.88 ;
      RECT 14.03 53.79 65.855 54.745 ;
      RECT 14.03 50.87 15.995 53.79 ;
      RECT 14.03 49.895 64.885 50.87 ;
      RECT 14.03 44.73 65.86 49.895 ;
      RECT 14.03 43.77 65.86 44.73 ;
      RECT 14.03 40.85 15.995 43.77 ;
      RECT 14.03 39.875 64.885 40.85 ;
      RECT 14.03 34.75 65.86 39.875 ;
      RECT 14.03 33.79 65.86 34.75 ;
      RECT 14.03 30.87 15.995 33.79 ;
      RECT 14.03 29.82 64.81 30.87 ;
      RECT 14.03 25.5 65.86 29.82 ;
      RECT 14.03 24.28 65.86 25.5 ;
      RECT 16.475 21.835 64.64 24.28 ;
      RECT 18.38 19.93 53.955 21.835 ;
      RECT 20.535 17.775 53.955 19.93 ;
      RECT 21.85 16.46 56.11 17.775 ;
      RECT 55.875 9.1 56.11 16.46 ;
      RECT 55.875 8.9 56.11 9.1 ;
      RECT 17.57 8.78 55.91 8.9 ;
      RECT 10.71 8.605 11.515 8.825 ;
      RECT 10.7 8.595 11.735 8.605 ;
      RECT 17.14 8.35 17.49 8.7 ;
      RECT 10.7 7.055 11.735 8.595 ;
      RECT 10.705 7.05 11.735 7.055 ;
      RECT 53.675 6.94 55.79 8.78 ;
      RECT 10.93 6.825 11.735 7.05 ;
      RECT 17.14 4.325 17.49 8.35 ;
      RECT 0 0 0.22 193.91 ;
      RECT 74.84 0 75 73.77 ;
      RECT 53.675 0 53.955 6.94 ;
      RECT 17.31 4.155 17.49 4.325 ;
      RECT 20.775 0.69 20.875 1.5 ;
      RECT 20.775 0 21.685 0.69 ;
      RECT 0 193.91 75 198 ;
      RECT 18.58 193.77 75 193.91 ;
      RECT 68.15 190.85 75 193.77 ;
      RECT 15.52 190.71 75 190.85 ;
      RECT 14.24 189.825 75 190.71 ;
      RECT 14.24 184.795 75 189.825 ;
      RECT 15.125 183.91 75 184.795 ;
      RECT 15.66 183.77 75 183.91 ;
      RECT 68.15 180.85 75 183.77 ;
      RECT 15.52 180.71 75 180.85 ;
      RECT 14.24 179.825 75 180.71 ;
      RECT 14.24 174.795 75 179.825 ;
      RECT 15.125 173.91 75 174.795 ;
      RECT 15.66 173.77 75 173.91 ;
      RECT 68.15 170.85 75 173.77 ;
      RECT 15.52 170.71 75 170.85 ;
      RECT 14.24 169.825 75 170.71 ;
      RECT 14.24 164.795 75 169.825 ;
      RECT 15.125 163.91 75 164.795 ;
      RECT 15.66 163.77 75 163.91 ;
      RECT 68.15 160.85 75 163.77 ;
      RECT 15.52 160.71 75 160.85 ;
      RECT 14.24 159.825 75 160.71 ;
      RECT 14.24 154.795 75 159.825 ;
      RECT 15.125 153.91 75 154.795 ;
      RECT 15.66 153.77 75 153.91 ;
      RECT 68.15 150.85 75 153.77 ;
      RECT 15.52 150.71 75 150.85 ;
      RECT 14.24 149.825 75 150.71 ;
      RECT 14.03 44.68 65.615 44.75 ;
      RECT 14.03 44.75 65.685 44.785 ;
      RECT 14.03 39.82 65.65 39.89 ;
      RECT 14.03 39.89 65.58 39.96 ;
      RECT 14.03 39.96 65.51 40.03 ;
      RECT 14.03 40.03 65.44 40.1 ;
      RECT 14.03 40.1 65.37 40.17 ;
      RECT 14.03 40.17 65.3 40.24 ;
      RECT 14.03 40.24 65.23 40.31 ;
      RECT 14.03 40.31 65.16 40.38 ;
      RECT 14.03 40.38 65.09 40.45 ;
      RECT 14.03 40.45 65.02 40.52 ;
      RECT 14.03 40.52 64.95 40.59 ;
      RECT 14.03 40.59 64.88 40.66 ;
      RECT 14.03 40.66 64.83 40.71 ;
      RECT 14.03 33.93 64.845 34 ;
      RECT 14.03 34 64.915 34.07 ;
      RECT 14.03 34.07 64.985 34.14 ;
      RECT 14.03 34.14 65.055 34.21 ;
      RECT 14.03 34.21 65.125 34.28 ;
      RECT 14.03 34.28 65.195 34.35 ;
      RECT 14.03 34.35 65.265 34.42 ;
      RECT 14.03 34.42 65.335 34.49 ;
      RECT 14.03 34.49 65.405 34.56 ;
      RECT 14.03 34.56 65.475 34.63 ;
      RECT 14.03 34.63 65.545 34.7 ;
      RECT 14.03 34.7 65.615 34.77 ;
      RECT 14.03 34.77 65.685 34.805 ;
      RECT 14.03 29.765 65.65 29.835 ;
      RECT 14.03 29.835 65.58 29.905 ;
      RECT 14.03 29.905 65.51 29.975 ;
      RECT 14.03 29.975 65.44 30.045 ;
      RECT 14.03 30.045 65.37 30.115 ;
      RECT 14.03 30.115 65.3 30.185 ;
      RECT 14.03 30.185 65.23 30.255 ;
      RECT 14.03 30.255 65.16 30.325 ;
      RECT 14.03 30.325 65.09 30.395 ;
      RECT 14.03 30.395 65.02 30.465 ;
      RECT 14.03 30.465 64.95 30.535 ;
      RECT 14.03 30.535 64.88 30.605 ;
      RECT 14.03 30.605 64.81 30.675 ;
      RECT 14.03 30.675 64.755 30.73 ;
      RECT 14.03 24.28 64.445 24.35 ;
      RECT 14.03 24.35 64.515 24.42 ;
      RECT 14.03 24.42 64.585 24.49 ;
      RECT 14.03 24.49 64.655 24.56 ;
      RECT 14.03 24.56 64.725 24.63 ;
      RECT 14.03 24.63 64.795 24.7 ;
      RECT 14.03 24.7 64.865 24.77 ;
      RECT 14.03 24.77 64.935 24.84 ;
      RECT 14.03 24.84 65.005 24.91 ;
      RECT 14.03 24.91 65.075 24.98 ;
      RECT 14.03 24.98 65.145 25.05 ;
      RECT 14.03 25.05 65.215 25.12 ;
      RECT 14.03 25.12 65.285 25.19 ;
      RECT 14.03 25.19 65.355 25.26 ;
      RECT 14.03 25.26 65.425 25.33 ;
      RECT 14.03 25.33 65.495 25.4 ;
      RECT 14.03 25.4 65.565 25.47 ;
      RECT 14.03 25.47 65.635 25.54 ;
      RECT 14.03 25.54 65.705 25.555 ;
      RECT 14.66 130.175 75 130.245 ;
      RECT 14.73 130.245 75 130.315 ;
      RECT 14.8 130.315 75 130.385 ;
      RECT 14.87 130.385 75 130.455 ;
      RECT 14.94 130.455 75 130.525 ;
      RECT 15.01 130.525 75 130.595 ;
      RECT 15.08 130.595 75 130.665 ;
      RECT 15.125 130.665 75 130.71 ;
      RECT 15.78 123.255 75 123.325 ;
      RECT 15.71 123.325 75 123.395 ;
      RECT 15.64 123.395 75 123.465 ;
      RECT 15.57 123.465 75 123.535 ;
      RECT 15.5 123.535 75 123.605 ;
      RECT 15.43 123.605 75 123.675 ;
      RECT 15.36 123.675 75 123.745 ;
      RECT 15.29 123.745 75 123.815 ;
      RECT 15.22 123.815 75 123.885 ;
      RECT 15.15 123.885 75 123.955 ;
      RECT 15.08 123.955 75 124.025 ;
      RECT 15.01 124.025 75 124.095 ;
      RECT 14.94 124.095 75 124.165 ;
      RECT 14.87 124.165 75 124.235 ;
      RECT 14.8 124.235 75 124.305 ;
      RECT 14.73 124.305 75 124.375 ;
      RECT 14.66 124.375 75 124.445 ;
      RECT 14.59 124.445 75 124.515 ;
      RECT 14.52 124.515 75 124.585 ;
      RECT 14.45 124.585 75 124.655 ;
      RECT 14.38 124.655 75 124.725 ;
      RECT 14.31 124.725 75 124.795 ;
      RECT 15.78 74.18 65.35 74.25 ;
      RECT 15.78 74.25 65.425 74.32 ;
      RECT 15.78 74.32 65.495 74.39 ;
      RECT 15.78 74.39 65.565 74.46 ;
      RECT 15.78 74.46 65.635 74.53 ;
      RECT 15.78 74.53 65.705 74.545 ;
      RECT 68.925 73.91 75 73.98 ;
      RECT 68.855 73.98 75 74.05 ;
      RECT 68.785 74.05 75 74.12 ;
      RECT 68.715 74.12 75 74.19 ;
      RECT 68.645 74.19 75 74.26 ;
      RECT 68.575 74.26 75 74.33 ;
      RECT 68.505 74.33 75 74.4 ;
      RECT 68.435 74.4 75 74.47 ;
      RECT 68.365 74.47 75 74.54 ;
      RECT 68.295 74.54 75 74.545 ;
      RECT 14.03 69.825 65.645 69.895 ;
      RECT 14.03 69.895 65.575 69.965 ;
      RECT 14.03 69.965 65.505 70.035 ;
      RECT 14.03 70.035 65.435 70.105 ;
      RECT 14.03 70.105 65.365 70.175 ;
      RECT 14.03 70.175 65.295 70.245 ;
      RECT 14.03 70.245 65.225 70.315 ;
      RECT 14.03 70.315 65.155 70.385 ;
      RECT 14.03 70.385 65.085 70.455 ;
      RECT 14.03 70.455 65.015 70.525 ;
      RECT 14.03 70.525 64.945 70.595 ;
      RECT 14.03 70.595 64.875 70.665 ;
      RECT 14.03 70.665 64.83 70.71 ;
      RECT 14.03 63.91 64.83 63.98 ;
      RECT 14.03 63.98 64.9 64.05 ;
      RECT 14.03 64.05 64.97 64.12 ;
      RECT 14.03 64.12 65.04 64.19 ;
      RECT 14.03 64.19 65.11 64.26 ;
      RECT 14.03 64.26 65.18 64.33 ;
      RECT 14.03 64.33 65.25 64.4 ;
      RECT 14.03 64.4 65.32 64.47 ;
      RECT 14.03 64.47 65.39 64.54 ;
      RECT 14.03 64.54 65.46 64.61 ;
      RECT 14.03 64.61 65.53 64.68 ;
      RECT 14.03 64.68 65.6 64.75 ;
      RECT 14.03 64.75 65.67 64.795 ;
      RECT 14.03 59.825 65.645 59.895 ;
      RECT 14.03 59.895 65.575 59.965 ;
      RECT 14.03 59.965 65.505 60.035 ;
      RECT 14.03 60.035 65.435 60.105 ;
      RECT 14.03 60.105 65.365 60.175 ;
      RECT 14.03 60.175 65.295 60.245 ;
      RECT 14.03 60.245 65.225 60.315 ;
      RECT 14.03 60.315 65.155 60.385 ;
      RECT 14.03 60.385 65.085 60.455 ;
      RECT 14.03 60.455 65.015 60.525 ;
      RECT 14.03 60.525 64.945 60.595 ;
      RECT 14.03 60.595 64.875 60.665 ;
      RECT 14.03 60.665 64.83 60.71 ;
      RECT 14.03 53.93 64.845 54 ;
      RECT 14.03 54 64.915 54.07 ;
      RECT 14.03 54.07 64.985 54.14 ;
      RECT 14.03 54.14 65.055 54.21 ;
      RECT 14.03 54.21 65.125 54.28 ;
      RECT 14.03 54.28 65.195 54.35 ;
      RECT 14.03 54.35 65.265 54.42 ;
      RECT 14.03 54.42 65.335 54.49 ;
      RECT 14.03 54.49 65.405 54.56 ;
      RECT 14.03 54.56 65.475 54.63 ;
      RECT 14.03 54.63 65.545 54.7 ;
      RECT 14.03 54.7 65.615 54.77 ;
      RECT 14.03 54.77 65.685 54.8 ;
      RECT 14.03 49.84 65.65 49.91 ;
      RECT 14.03 49.91 65.58 49.98 ;
      RECT 14.03 49.98 65.51 50.05 ;
      RECT 14.03 50.05 65.44 50.12 ;
      RECT 14.03 50.12 65.37 50.19 ;
      RECT 14.03 50.19 65.3 50.26 ;
      RECT 14.03 50.26 65.23 50.33 ;
      RECT 14.03 50.33 65.16 50.4 ;
      RECT 14.03 50.4 65.09 50.47 ;
      RECT 14.03 50.47 65.02 50.54 ;
      RECT 14.03 50.54 64.95 50.61 ;
      RECT 14.03 50.61 64.88 50.68 ;
      RECT 14.03 50.68 64.83 50.73 ;
      RECT 14.03 43.91 64.845 43.98 ;
      RECT 14.03 43.98 64.915 44.05 ;
      RECT 14.03 44.05 64.985 44.12 ;
      RECT 14.03 44.12 65.055 44.19 ;
      RECT 14.03 44.19 65.125 44.26 ;
      RECT 14.03 44.26 65.195 44.33 ;
      RECT 14.03 44.33 65.265 44.4 ;
      RECT 14.03 44.4 65.335 44.47 ;
      RECT 14.03 44.47 65.405 44.54 ;
      RECT 14.03 44.54 65.475 44.61 ;
      RECT 14.03 44.61 65.545 44.68 ;
      RECT 15.125 173.91 75 173.98 ;
      RECT 15.055 173.98 75 174.05 ;
      RECT 14.985 174.05 75 174.12 ;
      RECT 14.915 174.12 75 174.19 ;
      RECT 14.845 174.19 75 174.26 ;
      RECT 14.775 174.26 75 174.33 ;
      RECT 14.705 174.33 75 174.4 ;
      RECT 14.635 174.4 75 174.47 ;
      RECT 14.565 174.47 75 174.54 ;
      RECT 14.495 174.54 75 174.61 ;
      RECT 14.425 174.61 75 174.68 ;
      RECT 14.355 174.68 75 174.75 ;
      RECT 14.285 174.75 75 174.795 ;
      RECT 14.31 169.825 75 169.895 ;
      RECT 14.38 169.895 75 169.965 ;
      RECT 14.45 169.965 75 170.035 ;
      RECT 14.52 170.035 75 170.105 ;
      RECT 14.59 170.105 75 170.175 ;
      RECT 14.66 170.175 75 170.245 ;
      RECT 14.73 170.245 75 170.315 ;
      RECT 14.8 170.315 75 170.385 ;
      RECT 14.87 170.385 75 170.455 ;
      RECT 14.94 170.455 75 170.525 ;
      RECT 15.01 170.525 75 170.595 ;
      RECT 15.08 170.595 75 170.665 ;
      RECT 15.125 170.665 75 170.71 ;
      RECT 15.125 163.91 75 163.98 ;
      RECT 15.055 163.98 75 164.05 ;
      RECT 14.985 164.05 75 164.12 ;
      RECT 14.915 164.12 75 164.19 ;
      RECT 14.845 164.19 75 164.26 ;
      RECT 14.775 164.26 75 164.33 ;
      RECT 14.705 164.33 75 164.4 ;
      RECT 14.635 164.4 75 164.47 ;
      RECT 14.565 164.47 75 164.54 ;
      RECT 14.495 164.54 75 164.61 ;
      RECT 14.425 164.61 75 164.68 ;
      RECT 14.355 164.68 75 164.75 ;
      RECT 14.285 164.75 75 164.795 ;
      RECT 14.31 159.825 75 159.895 ;
      RECT 14.38 159.895 75 159.965 ;
      RECT 14.45 159.965 75 160.035 ;
      RECT 14.52 160.035 75 160.105 ;
      RECT 14.59 160.105 75 160.175 ;
      RECT 14.66 160.175 75 160.245 ;
      RECT 14.73 160.245 75 160.315 ;
      RECT 14.8 160.315 75 160.385 ;
      RECT 14.87 160.385 75 160.455 ;
      RECT 14.94 160.455 75 160.525 ;
      RECT 15.01 160.525 75 160.595 ;
      RECT 15.08 160.595 75 160.665 ;
      RECT 15.125 160.665 75 160.71 ;
      RECT 15.125 153.91 75 153.98 ;
      RECT 15.055 153.98 75 154.05 ;
      RECT 14.985 154.05 75 154.12 ;
      RECT 14.915 154.12 75 154.19 ;
      RECT 14.845 154.19 75 154.26 ;
      RECT 14.775 154.26 75 154.33 ;
      RECT 14.705 154.33 75 154.4 ;
      RECT 14.635 154.4 75 154.47 ;
      RECT 14.565 154.47 75 154.54 ;
      RECT 14.495 154.54 75 154.61 ;
      RECT 14.425 154.61 75 154.68 ;
      RECT 14.355 154.68 75 154.75 ;
      RECT 14.285 154.75 75 154.795 ;
      RECT 14.31 149.825 75 149.895 ;
      RECT 14.38 149.895 75 149.965 ;
      RECT 14.45 149.965 75 150.035 ;
      RECT 14.52 150.035 75 150.105 ;
      RECT 14.59 150.105 75 150.175 ;
      RECT 14.66 150.175 75 150.245 ;
      RECT 14.73 150.245 75 150.315 ;
      RECT 14.8 150.315 75 150.385 ;
      RECT 14.87 150.385 75 150.455 ;
      RECT 14.94 150.455 75 150.525 ;
      RECT 15.01 150.525 75 150.595 ;
      RECT 15.08 150.595 75 150.665 ;
      RECT 15.125 150.665 75 150.71 ;
      RECT 15.125 143.91 75 143.98 ;
      RECT 15.055 143.98 75 144.05 ;
      RECT 14.985 144.05 75 144.12 ;
      RECT 14.915 144.12 75 144.19 ;
      RECT 14.845 144.19 75 144.26 ;
      RECT 14.775 144.26 75 144.33 ;
      RECT 14.705 144.33 75 144.4 ;
      RECT 14.635 144.4 75 144.47 ;
      RECT 14.565 144.47 75 144.54 ;
      RECT 14.495 144.54 75 144.61 ;
      RECT 14.425 144.61 75 144.68 ;
      RECT 14.355 144.68 75 144.75 ;
      RECT 14.285 144.75 75 144.795 ;
      RECT 14.31 139.825 75 139.895 ;
      RECT 14.38 139.895 75 139.965 ;
      RECT 14.45 139.965 75 140.035 ;
      RECT 14.52 140.035 75 140.105 ;
      RECT 14.59 140.105 75 140.175 ;
      RECT 14.66 140.175 75 140.245 ;
      RECT 14.73 140.245 75 140.315 ;
      RECT 14.8 140.315 75 140.385 ;
      RECT 14.87 140.385 75 140.455 ;
      RECT 14.94 140.455 75 140.525 ;
      RECT 15.01 140.525 75 140.595 ;
      RECT 15.08 140.595 75 140.665 ;
      RECT 15.125 140.665 75 140.71 ;
      RECT 15.125 133.91 75 133.98 ;
      RECT 15.055 133.98 75 134.05 ;
      RECT 14.985 134.05 75 134.12 ;
      RECT 14.915 134.12 75 134.19 ;
      RECT 14.845 134.19 75 134.26 ;
      RECT 14.775 134.26 75 134.33 ;
      RECT 14.705 134.33 75 134.4 ;
      RECT 14.635 134.4 75 134.47 ;
      RECT 14.565 134.47 75 134.54 ;
      RECT 14.495 134.54 75 134.61 ;
      RECT 14.425 134.61 75 134.68 ;
      RECT 14.355 134.68 75 134.75 ;
      RECT 14.285 134.75 75 134.795 ;
      RECT 14.31 129.825 75 129.895 ;
      RECT 14.38 129.895 75 129.965 ;
      RECT 14.45 129.965 75 130.035 ;
      RECT 14.52 130.035 75 130.105 ;
      RECT 14.59 130.105 75 130.175 ;
      RECT 16.125 22.185 62.35 22.255 ;
      RECT 16.195 22.115 62.28 22.185 ;
      RECT 16.265 22.045 62.21 22.115 ;
      RECT 16.335 21.975 62.14 22.045 ;
      RECT 18.435 19.875 53.815 19.945 ;
      RECT 18.365 19.945 53.815 20.015 ;
      RECT 18.295 20.015 53.815 20.085 ;
      RECT 18.225 20.085 53.815 20.155 ;
      RECT 18.155 20.155 53.815 20.225 ;
      RECT 18.085 20.225 53.815 20.295 ;
      RECT 18.015 20.295 53.815 20.365 ;
      RECT 17.945 20.365 53.815 20.435 ;
      RECT 17.875 20.435 53.815 20.505 ;
      RECT 17.805 20.505 53.815 20.575 ;
      RECT 17.735 20.575 53.815 20.645 ;
      RECT 17.665 20.645 53.815 20.715 ;
      RECT 17.595 20.715 53.815 20.785 ;
      RECT 17.525 20.785 53.815 20.855 ;
      RECT 17.455 20.855 53.815 20.925 ;
      RECT 17.385 20.925 53.815 20.995 ;
      RECT 17.315 20.995 53.815 21.065 ;
      RECT 17.245 21.065 53.815 21.135 ;
      RECT 17.175 21.135 53.815 21.205 ;
      RECT 17.105 21.205 53.815 21.275 ;
      RECT 17.035 21.275 53.815 21.345 ;
      RECT 16.965 21.345 53.815 21.415 ;
      RECT 16.895 21.415 53.815 21.485 ;
      RECT 16.825 21.485 53.815 21.555 ;
      RECT 16.755 21.555 53.815 21.625 ;
      RECT 16.685 21.625 53.815 21.695 ;
      RECT 16.615 21.695 53.815 21.765 ;
      RECT 16.545 21.765 53.815 21.835 ;
      RECT 16.475 21.835 53.815 21.905 ;
      RECT 16.405 21.905 53.815 21.975 ;
      RECT 20.59 17.72 55.9 17.79 ;
      RECT 20.52 17.79 55.83 17.86 ;
      RECT 20.45 17.86 55.76 17.93 ;
      RECT 20.38 17.93 55.69 18 ;
      RECT 20.31 18 55.62 18.07 ;
      RECT 20.24 18.07 55.55 18.14 ;
      RECT 20.17 18.14 55.48 18.21 ;
      RECT 20.1 18.21 55.41 18.28 ;
      RECT 20.03 18.28 55.34 18.35 ;
      RECT 19.96 18.35 55.27 18.42 ;
      RECT 19.89 18.42 55.2 18.49 ;
      RECT 19.82 18.49 55.13 18.56 ;
      RECT 19.75 18.56 55.06 18.63 ;
      RECT 19.68 18.63 54.99 18.7 ;
      RECT 19.61 18.7 54.92 18.77 ;
      RECT 19.54 18.77 54.85 18.84 ;
      RECT 19.47 18.84 54.78 18.91 ;
      RECT 19.4 18.91 54.71 18.98 ;
      RECT 19.33 18.98 54.64 19.05 ;
      RECT 19.26 19.05 54.57 19.12 ;
      RECT 19.19 19.12 54.5 19.19 ;
      RECT 19.12 19.19 54.43 19.26 ;
      RECT 19.05 19.26 54.36 19.33 ;
      RECT 18.98 19.33 54.29 19.4 ;
      RECT 18.91 19.4 54.22 19.47 ;
      RECT 18.84 19.47 54.15 19.54 ;
      RECT 18.77 19.54 54.08 19.61 ;
      RECT 18.7 19.61 54.01 19.68 ;
      RECT 18.63 19.68 53.94 19.75 ;
      RECT 18.56 19.75 53.87 19.82 ;
      RECT 18.49 19.82 53.815 19.875 ;
      RECT 21.85 16.46 55.97 16.53 ;
      RECT 21.78 16.53 55.97 16.6 ;
      RECT 21.71 16.6 55.97 16.67 ;
      RECT 21.64 16.67 55.97 16.74 ;
      RECT 21.57 16.74 55.97 16.81 ;
      RECT 21.5 16.81 55.97 16.88 ;
      RECT 21.43 16.88 55.97 16.95 ;
      RECT 21.36 16.95 55.97 17.02 ;
      RECT 21.29 17.02 55.97 17.09 ;
      RECT 21.22 17.09 55.97 17.16 ;
      RECT 21.15 17.16 55.97 17.23 ;
      RECT 21.08 17.23 55.97 17.3 ;
      RECT 21.01 17.3 55.97 17.37 ;
      RECT 20.94 17.37 55.97 17.44 ;
      RECT 20.87 17.44 55.97 17.51 ;
      RECT 20.8 17.51 55.97 17.58 ;
      RECT 20.73 17.58 55.97 17.65 ;
      RECT 20.66 17.65 55.97 17.72 ;
      RECT 15.78 73.91 65.085 73.98 ;
      RECT 15.78 73.98 65.155 74.05 ;
      RECT 15.78 74.05 65.225 74.12 ;
      RECT 15.78 74.12 65.295 74.18 ;
      RECT 14.31 189.825 75 189.895 ;
      RECT 14.38 189.895 75 189.965 ;
      RECT 14.45 189.965 75 190.035 ;
      RECT 14.52 190.035 75 190.105 ;
      RECT 14.59 190.105 75 190.175 ;
      RECT 14.66 190.175 75 190.245 ;
      RECT 14.73 190.245 75 190.315 ;
      RECT 14.8 190.315 75 190.385 ;
      RECT 14.87 190.385 75 190.455 ;
      RECT 14.94 190.455 75 190.525 ;
      RECT 15.01 190.525 75 190.595 ;
      RECT 15.08 190.595 75 190.665 ;
      RECT 15.125 190.665 75 190.71 ;
      RECT 15.125 183.91 75 183.98 ;
      RECT 15.055 183.98 75 184.05 ;
      RECT 14.985 184.05 75 184.12 ;
      RECT 14.915 184.12 75 184.19 ;
      RECT 14.845 184.19 75 184.26 ;
      RECT 14.775 184.26 75 184.33 ;
      RECT 14.705 184.33 75 184.4 ;
      RECT 14.635 184.4 75 184.47 ;
      RECT 14.565 184.47 75 184.54 ;
      RECT 14.495 184.54 75 184.61 ;
      RECT 14.425 184.61 75 184.68 ;
      RECT 14.355 184.68 75 184.75 ;
      RECT 14.285 184.75 75 184.795 ;
      RECT 14.31 179.825 75 179.895 ;
      RECT 14.38 179.895 75 179.965 ;
      RECT 14.45 179.965 75 180.035 ;
      RECT 14.52 180.035 75 180.105 ;
      RECT 14.59 180.105 75 180.175 ;
      RECT 14.66 180.175 75 180.245 ;
      RECT 14.73 180.245 75 180.315 ;
      RECT 14.8 180.315 75 180.385 ;
      RECT 14.87 180.385 75 180.455 ;
      RECT 14.94 180.455 75 180.525 ;
      RECT 15.01 180.525 75 180.595 ;
      RECT 15.08 180.595 75 180.665 ;
      RECT 15.125 180.665 75 180.71 ;
      RECT 15.145 23.165 63.33 23.235 ;
      RECT 15.215 23.095 63.26 23.165 ;
      RECT 15.285 23.025 63.19 23.095 ;
      RECT 15.355 22.955 63.12 23.025 ;
      RECT 15.425 22.885 63.05 22.955 ;
      RECT 15.495 22.815 62.98 22.885 ;
      RECT 15.565 22.745 62.91 22.815 ;
      RECT 15.635 22.675 62.84 22.745 ;
      RECT 15.705 22.605 62.77 22.675 ;
      RECT 15.775 22.535 62.7 22.605 ;
      RECT 15.845 22.465 62.63 22.535 ;
      RECT 15.915 22.395 62.56 22.465 ;
      RECT 15.985 22.325 62.49 22.395 ;
      RECT 16.055 22.255 62.42 22.325 ;
      RECT 16.125 22.185 62.35 22.255 ;
      RECT 16.195 22.115 62.28 22.185 ;
      RECT 16.265 22.045 62.21 22.115 ;
      RECT 16.335 21.975 62.14 22.045 ;
      RECT 18.435 19.875 53.815 19.945 ;
      RECT 18.365 19.945 53.815 20.015 ;
      RECT 18.295 20.015 53.815 20.085 ;
      RECT 18.225 20.085 53.815 20.155 ;
      RECT 18.155 20.155 53.815 20.225 ;
      RECT 18.085 20.225 53.815 20.295 ;
      RECT 18.015 20.295 53.815 20.365 ;
      RECT 17.945 20.365 53.815 20.435 ;
      RECT 17.875 20.435 53.815 20.505 ;
      RECT 17.805 20.505 53.815 20.575 ;
      RECT 17.735 20.575 53.815 20.645 ;
      RECT 17.665 20.645 53.815 20.715 ;
      RECT 17.595 20.715 53.815 20.785 ;
      RECT 17.525 20.785 53.815 20.855 ;
      RECT 17.455 20.855 53.815 20.925 ;
      RECT 17.385 20.925 53.815 20.995 ;
      RECT 17.315 20.995 53.815 21.065 ;
      RECT 17.245 21.065 53.815 21.135 ;
      RECT 17.175 21.135 53.815 21.205 ;
      RECT 17.105 21.205 53.815 21.275 ;
      RECT 17.035 21.275 53.815 21.345 ;
      RECT 16.965 21.345 53.815 21.415 ;
      RECT 16.895 21.415 53.815 21.485 ;
      RECT 16.825 21.485 53.815 21.555 ;
      RECT 16.755 21.555 53.815 21.625 ;
      RECT 16.685 21.625 53.815 21.695 ;
      RECT 16.615 21.695 53.815 21.765 ;
      RECT 16.545 21.765 53.815 21.835 ;
      RECT 16.475 21.835 53.815 21.905 ;
      RECT 16.405 21.905 53.815 21.975 ;
      RECT 20.59 17.72 55.9 17.79 ;
      RECT 20.52 17.79 55.83 17.86 ;
      RECT 20.45 17.86 55.76 17.93 ;
      RECT 20.38 17.93 55.69 18 ;
      RECT 20.31 18 55.62 18.07 ;
      RECT 20.24 18.07 55.55 18.14 ;
      RECT 20.17 18.14 55.48 18.21 ;
      RECT 20.1 18.21 55.41 18.28 ;
      RECT 20.03 18.28 55.34 18.35 ;
      RECT 19.96 18.35 55.27 18.42 ;
      RECT 19.89 18.42 55.2 18.49 ;
      RECT 19.82 18.49 55.13 18.56 ;
      RECT 19.75 18.56 55.06 18.63 ;
      RECT 19.68 18.63 54.99 18.7 ;
      RECT 19.61 18.7 54.92 18.77 ;
      RECT 19.54 18.77 54.85 18.84 ;
      RECT 19.47 18.84 54.78 18.91 ;
      RECT 19.4 18.91 54.71 18.98 ;
      RECT 19.33 18.98 54.64 19.05 ;
      RECT 19.26 19.05 54.57 19.12 ;
      RECT 19.19 19.12 54.5 19.19 ;
      RECT 19.12 19.19 54.43 19.26 ;
      RECT 19.05 19.26 54.36 19.33 ;
      RECT 18.98 19.33 54.29 19.4 ;
      RECT 18.91 19.4 54.22 19.47 ;
      RECT 18.84 19.47 54.15 19.54 ;
      RECT 18.77 19.54 54.08 19.61 ;
      RECT 18.7 19.61 54.01 19.68 ;
      RECT 18.63 19.68 53.94 19.75 ;
      RECT 18.56 19.75 53.87 19.82 ;
      RECT 18.49 19.82 53.815 19.875 ;
      RECT 21.85 16.46 55.97 16.53 ;
      RECT 21.78 16.53 55.97 16.6 ;
      RECT 21.71 16.6 55.97 16.67 ;
      RECT 21.64 16.67 55.97 16.74 ;
      RECT 21.57 16.74 55.97 16.81 ;
      RECT 21.5 16.81 55.97 16.88 ;
      RECT 21.43 16.88 55.97 16.95 ;
      RECT 21.36 16.95 55.97 17.02 ;
      RECT 21.29 17.02 55.97 17.09 ;
      RECT 21.22 17.09 55.97 17.16 ;
      RECT 21.15 17.16 55.97 17.23 ;
      RECT 21.08 17.23 55.97 17.3 ;
      RECT 21.01 17.3 55.97 17.37 ;
      RECT 20.94 17.37 55.97 17.44 ;
      RECT 20.87 17.44 55.97 17.51 ;
      RECT 20.8 17.51 55.97 17.58 ;
      RECT 20.73 17.58 55.97 17.65 ;
      RECT 20.66 17.65 55.97 17.72 ;
      RECT 14.095 24.215 64.38 24.28 ;
      RECT 14.165 24.145 64.31 24.215 ;
      RECT 14.235 24.075 64.24 24.145 ;
      RECT 14.305 24.005 64.17 24.075 ;
      RECT 14.375 23.935 64.1 24.005 ;
      RECT 14.445 23.865 64.03 23.935 ;
      RECT 14.515 23.795 63.96 23.865 ;
      RECT 14.585 23.725 63.89 23.795 ;
      RECT 14.655 23.655 63.82 23.725 ;
      RECT 14.725 23.585 63.75 23.655 ;
      RECT 14.795 23.515 63.68 23.585 ;
      RECT 14.865 23.445 63.61 23.515 ;
      RECT 14.935 23.375 63.54 23.445 ;
      RECT 15.005 23.305 63.47 23.375 ;
      RECT 15.075 23.235 63.4 23.305 ;
      RECT 15.145 23.165 63.33 23.235 ;
      RECT 15.215 23.095 63.26 23.165 ;
      RECT 15.285 23.025 63.19 23.095 ;
      RECT 15.355 22.955 63.12 23.025 ;
      RECT 15.425 22.885 63.05 22.955 ;
      RECT 15.495 22.815 62.98 22.885 ;
      RECT 15.565 22.745 62.91 22.815 ;
      RECT 15.635 22.675 62.84 22.745 ;
      RECT 15.705 22.605 62.77 22.675 ;
      RECT 15.775 22.535 62.7 22.605 ;
      RECT 15.845 22.465 62.63 22.535 ;
      RECT 15.915 22.395 62.56 22.465 ;
      RECT 15.985 22.325 62.49 22.395 ;
      RECT 16.055 22.255 62.42 22.325 ;
      RECT 14.03 60.105 65.365 60.175 ;
      RECT 14.03 60.175 65.295 60.245 ;
      RECT 14.03 60.245 65.225 60.315 ;
      RECT 14.03 60.315 65.155 60.385 ;
      RECT 14.03 60.385 65.085 60.455 ;
      RECT 14.03 60.455 65.015 60.525 ;
      RECT 14.03 60.525 64.945 60.595 ;
      RECT 14.03 60.595 64.875 60.665 ;
      RECT 14.03 60.665 64.83 60.71 ;
      RECT 14.03 53.93 64.845 54 ;
      RECT 14.03 54 64.915 54.07 ;
      RECT 14.03 54.07 64.985 54.14 ;
      RECT 14.03 54.14 65.055 54.21 ;
      RECT 14.03 54.21 65.125 54.28 ;
      RECT 14.03 54.28 65.195 54.35 ;
      RECT 14.03 54.35 65.265 54.42 ;
      RECT 14.03 54.42 65.335 54.49 ;
      RECT 14.03 54.49 65.405 54.56 ;
      RECT 14.03 54.56 65.475 54.63 ;
      RECT 14.03 54.63 65.545 54.7 ;
      RECT 14.03 54.7 65.615 54.77 ;
      RECT 14.03 54.77 65.685 54.8 ;
      RECT 14.03 49.84 65.65 49.91 ;
      RECT 14.03 49.91 65.58 49.98 ;
      RECT 14.03 49.98 65.51 50.05 ;
      RECT 14.03 50.05 65.44 50.12 ;
      RECT 14.03 50.12 65.37 50.19 ;
      RECT 14.03 50.19 65.3 50.26 ;
      RECT 14.03 50.26 65.23 50.33 ;
      RECT 14.03 50.33 65.16 50.4 ;
      RECT 14.03 50.4 65.09 50.47 ;
      RECT 14.03 50.47 65.02 50.54 ;
      RECT 14.03 50.54 64.95 50.61 ;
      RECT 14.03 50.61 64.88 50.68 ;
      RECT 14.03 50.68 64.83 50.73 ;
      RECT 14.03 43.91 64.845 43.98 ;
      RECT 14.03 43.98 64.915 44.05 ;
      RECT 14.03 44.05 64.985 44.12 ;
      RECT 14.03 44.12 65.055 44.19 ;
      RECT 14.03 44.19 65.125 44.26 ;
      RECT 14.03 44.26 65.195 44.33 ;
      RECT 14.03 44.33 65.265 44.4 ;
      RECT 14.03 44.4 65.335 44.47 ;
      RECT 14.03 44.47 65.405 44.54 ;
      RECT 14.03 44.54 65.475 44.61 ;
      RECT 14.03 44.61 65.545 44.68 ;
      RECT 14.03 44.68 65.615 44.75 ;
      RECT 14.03 44.75 65.685 44.785 ;
      RECT 14.03 39.82 65.65 39.89 ;
      RECT 14.03 39.89 65.58 39.96 ;
      RECT 14.03 39.96 65.51 40.03 ;
      RECT 14.03 40.03 65.44 40.1 ;
      RECT 14.03 40.1 65.37 40.17 ;
      RECT 14.03 40.17 65.3 40.24 ;
      RECT 14.03 40.24 65.23 40.31 ;
      RECT 14.03 40.31 65.16 40.38 ;
      RECT 14.03 40.38 65.09 40.45 ;
      RECT 14.03 40.45 65.02 40.52 ;
      RECT 14.03 40.52 64.95 40.59 ;
      RECT 14.03 40.59 64.88 40.66 ;
      RECT 14.03 40.66 64.83 40.71 ;
      RECT 14.03 33.93 64.845 34 ;
      RECT 14.03 34 64.915 34.07 ;
      RECT 14.03 34.07 64.985 34.14 ;
      RECT 14.03 34.14 65.055 34.21 ;
      RECT 14.03 34.21 65.125 34.28 ;
      RECT 14.03 34.28 65.195 34.35 ;
      RECT 14.03 34.35 65.265 34.42 ;
      RECT 14.03 34.42 65.335 34.49 ;
      RECT 14.03 34.49 65.405 34.56 ;
      RECT 14.03 34.56 65.475 34.63 ;
      RECT 14.03 34.63 65.545 34.7 ;
      RECT 14.03 34.7 65.615 34.77 ;
      RECT 14.03 34.77 65.685 34.805 ;
      RECT 14.03 29.765 65.65 29.835 ;
      RECT 14.03 29.835 65.58 29.905 ;
      RECT 14.03 29.905 65.51 29.975 ;
      RECT 14.03 29.975 65.44 30.045 ;
      RECT 14.03 30.045 65.37 30.115 ;
      RECT 14.03 30.115 65.3 30.185 ;
      RECT 14.03 30.185 65.23 30.255 ;
      RECT 14.03 30.255 65.16 30.325 ;
      RECT 14.03 30.325 65.09 30.395 ;
      RECT 14.03 30.395 65.02 30.465 ;
      RECT 14.03 30.465 64.95 30.535 ;
      RECT 14.03 30.535 64.88 30.605 ;
      RECT 14.03 30.605 64.81 30.675 ;
      RECT 14.03 30.675 64.755 30.73 ;
      RECT 14.03 24.28 64.445 24.35 ;
      RECT 14.03 24.35 64.515 24.42 ;
      RECT 14.03 24.42 64.585 24.49 ;
      RECT 14.03 24.49 64.655 24.56 ;
      RECT 14.03 24.56 64.725 24.63 ;
      RECT 14.03 24.63 64.795 24.7 ;
      RECT 14.03 24.7 64.865 24.77 ;
      RECT 14.03 24.77 64.935 24.84 ;
      RECT 14.03 24.84 65.005 24.91 ;
      RECT 14.03 24.91 65.075 24.98 ;
      RECT 14.03 24.98 65.145 25.05 ;
      RECT 14.03 25.05 65.215 25.12 ;
      RECT 14.03 25.12 65.285 25.19 ;
      RECT 14.03 25.19 65.355 25.26 ;
      RECT 14.03 25.26 65.425 25.33 ;
      RECT 14.03 25.33 65.495 25.4 ;
      RECT 14.03 25.4 65.565 25.47 ;
      RECT 14.03 25.47 65.635 25.54 ;
      RECT 14.03 25.54 65.705 25.555 ;
      RECT 14.095 24.215 64.38 24.28 ;
      RECT 14.165 24.145 64.31 24.215 ;
      RECT 14.235 24.075 64.24 24.145 ;
      RECT 14.305 24.005 64.17 24.075 ;
      RECT 14.375 23.935 64.1 24.005 ;
      RECT 14.445 23.865 64.03 23.935 ;
      RECT 14.515 23.795 63.96 23.865 ;
      RECT 14.585 23.725 63.89 23.795 ;
      RECT 14.655 23.655 63.82 23.725 ;
      RECT 14.725 23.585 63.75 23.655 ;
      RECT 14.795 23.515 63.68 23.585 ;
      RECT 14.865 23.445 63.61 23.515 ;
      RECT 14.935 23.375 63.54 23.445 ;
      RECT 15.005 23.305 63.47 23.375 ;
      RECT 15.075 23.235 63.4 23.305 ;
      RECT 14.915 144.12 75 144.19 ;
      RECT 14.845 144.19 75 144.26 ;
      RECT 14.775 144.26 75 144.33 ;
      RECT 14.705 144.33 75 144.4 ;
      RECT 14.635 144.4 75 144.47 ;
      RECT 14.565 144.47 75 144.54 ;
      RECT 14.495 144.54 75 144.61 ;
      RECT 14.425 144.61 75 144.68 ;
      RECT 14.355 144.68 75 144.75 ;
      RECT 14.285 144.75 75 144.795 ;
      RECT 14.31 139.825 75 139.895 ;
      RECT 14.38 139.895 75 139.965 ;
      RECT 14.45 139.965 75 140.035 ;
      RECT 14.52 140.035 75 140.105 ;
      RECT 14.59 140.105 75 140.175 ;
      RECT 14.66 140.175 75 140.245 ;
      RECT 14.73 140.245 75 140.315 ;
      RECT 14.8 140.315 75 140.385 ;
      RECT 14.87 140.385 75 140.455 ;
      RECT 14.94 140.455 75 140.525 ;
      RECT 15.01 140.525 75 140.595 ;
      RECT 15.08 140.595 75 140.665 ;
      RECT 15.125 140.665 75 140.71 ;
      RECT 15.125 133.91 75 133.98 ;
      RECT 15.055 133.98 75 134.05 ;
      RECT 14.985 134.05 75 134.12 ;
      RECT 14.915 134.12 75 134.19 ;
      RECT 14.845 134.19 75 134.26 ;
      RECT 14.775 134.26 75 134.33 ;
      RECT 14.705 134.33 75 134.4 ;
      RECT 14.635 134.4 75 134.47 ;
      RECT 14.565 134.47 75 134.54 ;
      RECT 14.495 134.54 75 134.61 ;
      RECT 14.425 134.61 75 134.68 ;
      RECT 14.355 134.68 75 134.75 ;
      RECT 14.285 134.75 75 134.795 ;
      RECT 14.31 129.825 75 129.895 ;
      RECT 14.38 129.895 75 129.965 ;
      RECT 14.45 129.965 75 130.035 ;
      RECT 14.52 130.035 75 130.105 ;
      RECT 14.59 130.105 75 130.175 ;
      RECT 14.66 130.175 75 130.245 ;
      RECT 14.73 130.245 75 130.315 ;
      RECT 14.8 130.315 75 130.385 ;
      RECT 14.87 130.385 75 130.455 ;
      RECT 14.94 130.455 75 130.525 ;
      RECT 15.01 130.525 75 130.595 ;
      RECT 15.08 130.595 75 130.665 ;
      RECT 15.125 130.665 75 130.71 ;
      RECT 15.78 123.255 75 123.325 ;
      RECT 15.71 123.325 75 123.395 ;
      RECT 15.64 123.395 75 123.465 ;
      RECT 15.57 123.465 75 123.535 ;
      RECT 15.5 123.535 75 123.605 ;
      RECT 15.43 123.605 75 123.675 ;
      RECT 15.36 123.675 75 123.745 ;
      RECT 15.29 123.745 75 123.815 ;
      RECT 15.22 123.815 75 123.885 ;
      RECT 15.15 123.885 75 123.955 ;
      RECT 15.08 123.955 75 124.025 ;
      RECT 15.01 124.025 75 124.095 ;
      RECT 14.94 124.095 75 124.165 ;
      RECT 14.87 124.165 75 124.235 ;
      RECT 14.8 124.235 75 124.305 ;
      RECT 14.73 124.305 75 124.375 ;
      RECT 14.66 124.375 75 124.445 ;
      RECT 14.59 124.445 75 124.515 ;
      RECT 14.52 124.515 75 124.585 ;
      RECT 14.45 124.585 75 124.655 ;
      RECT 14.38 124.655 75 124.725 ;
      RECT 14.31 124.725 75 124.795 ;
      RECT 15.78 74.18 65.35 74.25 ;
      RECT 15.78 74.25 65.425 74.32 ;
      RECT 15.78 74.32 65.495 74.39 ;
      RECT 15.78 74.39 65.565 74.46 ;
      RECT 15.78 74.46 65.635 74.53 ;
      RECT 15.78 74.53 65.705 74.545 ;
      RECT 15.78 73.91 65.085 73.98 ;
      RECT 15.78 73.98 65.155 74.05 ;
      RECT 15.78 74.05 65.225 74.12 ;
      RECT 15.78 74.12 65.295 74.18 ;
      RECT 68.925 73.91 75 73.98 ;
      RECT 68.855 73.98 75 74.05 ;
      RECT 68.785 74.05 75 74.12 ;
      RECT 68.715 74.12 75 74.19 ;
      RECT 68.645 74.19 75 74.26 ;
      RECT 68.575 74.26 75 74.33 ;
      RECT 68.505 74.33 75 74.4 ;
      RECT 68.435 74.4 75 74.47 ;
      RECT 68.365 74.47 75 74.54 ;
      RECT 68.295 74.54 75 74.545 ;
      RECT 14.03 69.825 65.645 69.895 ;
      RECT 14.03 69.895 65.575 69.965 ;
      RECT 14.03 69.965 65.505 70.035 ;
      RECT 14.03 70.035 65.435 70.105 ;
      RECT 14.03 70.105 65.365 70.175 ;
      RECT 14.03 70.175 65.295 70.245 ;
      RECT 14.03 70.245 65.225 70.315 ;
      RECT 14.03 70.315 65.155 70.385 ;
      RECT 14.03 70.385 65.085 70.455 ;
      RECT 14.03 70.455 65.015 70.525 ;
      RECT 14.03 70.525 64.945 70.595 ;
      RECT 14.03 70.595 64.875 70.665 ;
      RECT 14.03 70.665 64.83 70.71 ;
      RECT 14.03 63.91 64.83 63.98 ;
      RECT 14.03 63.98 64.9 64.05 ;
      RECT 14.03 64.05 64.97 64.12 ;
      RECT 14.03 64.12 65.04 64.19 ;
      RECT 14.03 64.19 65.11 64.26 ;
      RECT 14.03 64.26 65.18 64.33 ;
      RECT 14.03 64.33 65.25 64.4 ;
      RECT 14.03 64.4 65.32 64.47 ;
      RECT 14.03 64.47 65.39 64.54 ;
      RECT 14.03 64.54 65.46 64.61 ;
      RECT 14.03 64.61 65.53 64.68 ;
      RECT 14.03 64.68 65.6 64.75 ;
      RECT 14.03 64.75 65.67 64.795 ;
      RECT 14.03 59.825 65.645 59.895 ;
      RECT 14.03 59.895 65.575 59.965 ;
      RECT 14.03 59.965 65.505 60.035 ;
      RECT 14.03 60.035 65.435 60.105 ;
      RECT 53.815 8.75 55.565 8.82 ;
      RECT 53.815 8.82 55.635 8.89 ;
      RECT 53.815 8.89 55.705 8.9 ;
      RECT 14.31 189.825 75 189.895 ;
      RECT 14.38 189.895 75 189.965 ;
      RECT 14.45 189.965 75 190.035 ;
      RECT 14.52 190.035 75 190.105 ;
      RECT 14.59 190.105 75 190.175 ;
      RECT 14.66 190.175 75 190.245 ;
      RECT 14.73 190.245 75 190.315 ;
      RECT 14.8 190.315 75 190.385 ;
      RECT 14.87 190.385 75 190.455 ;
      RECT 14.94 190.455 75 190.525 ;
      RECT 15.01 190.525 75 190.595 ;
      RECT 15.08 190.595 75 190.665 ;
      RECT 15.125 190.665 75 190.71 ;
      RECT 15.125 183.91 75 183.98 ;
      RECT 15.055 183.98 75 184.05 ;
      RECT 14.985 184.05 75 184.12 ;
      RECT 14.915 184.12 75 184.19 ;
      RECT 14.845 184.19 75 184.26 ;
      RECT 14.775 184.26 75 184.33 ;
      RECT 14.705 184.33 75 184.4 ;
      RECT 14.635 184.4 75 184.47 ;
      RECT 14.565 184.47 75 184.54 ;
      RECT 14.495 184.54 75 184.61 ;
      RECT 14.425 184.61 75 184.68 ;
      RECT 14.355 184.68 75 184.75 ;
      RECT 14.285 184.75 75 184.795 ;
      RECT 14.31 179.825 75 179.895 ;
      RECT 14.38 179.895 75 179.965 ;
      RECT 14.45 179.965 75 180.035 ;
      RECT 14.52 180.035 75 180.105 ;
      RECT 14.59 180.105 75 180.175 ;
      RECT 14.66 180.175 75 180.245 ;
      RECT 14.73 180.245 75 180.315 ;
      RECT 14.8 180.315 75 180.385 ;
      RECT 14.87 180.385 75 180.455 ;
      RECT 14.94 180.455 75 180.525 ;
      RECT 15.01 180.525 75 180.595 ;
      RECT 15.08 180.595 75 180.665 ;
      RECT 15.125 180.665 75 180.71 ;
      RECT 15.125 173.91 75 173.98 ;
      RECT 15.055 173.98 75 174.05 ;
      RECT 14.985 174.05 75 174.12 ;
      RECT 14.915 174.12 75 174.19 ;
      RECT 14.845 174.19 75 174.26 ;
      RECT 14.775 174.26 75 174.33 ;
      RECT 14.705 174.33 75 174.4 ;
      RECT 14.635 174.4 75 174.47 ;
      RECT 14.565 174.47 75 174.54 ;
      RECT 14.495 174.54 75 174.61 ;
      RECT 14.425 174.61 75 174.68 ;
      RECT 14.355 174.68 75 174.75 ;
      RECT 14.285 174.75 75 174.795 ;
      RECT 14.31 169.825 75 169.895 ;
      RECT 14.38 169.895 75 169.965 ;
      RECT 14.45 169.965 75 170.035 ;
      RECT 14.52 170.035 75 170.105 ;
      RECT 14.59 170.105 75 170.175 ;
      RECT 14.66 170.175 75 170.245 ;
      RECT 14.73 170.245 75 170.315 ;
      RECT 14.8 170.315 75 170.385 ;
      RECT 14.87 170.385 75 170.455 ;
      RECT 14.94 170.455 75 170.525 ;
      RECT 15.01 170.525 75 170.595 ;
      RECT 15.08 170.595 75 170.665 ;
      RECT 15.125 170.665 75 170.71 ;
      RECT 15.125 163.91 75 163.98 ;
      RECT 15.055 163.98 75 164.05 ;
      RECT 14.985 164.05 75 164.12 ;
      RECT 14.915 164.12 75 164.19 ;
      RECT 14.845 164.19 75 164.26 ;
      RECT 14.775 164.26 75 164.33 ;
      RECT 14.705 164.33 75 164.4 ;
      RECT 14.635 164.4 75 164.47 ;
      RECT 14.565 164.47 75 164.54 ;
      RECT 14.495 164.54 75 164.61 ;
      RECT 14.425 164.61 75 164.68 ;
      RECT 14.355 164.68 75 164.75 ;
      RECT 14.285 164.75 75 164.795 ;
      RECT 14.31 159.825 75 159.895 ;
      RECT 14.38 159.895 75 159.965 ;
      RECT 14.45 159.965 75 160.035 ;
      RECT 14.52 160.035 75 160.105 ;
      RECT 14.59 160.105 75 160.175 ;
      RECT 14.66 160.175 75 160.245 ;
      RECT 14.73 160.245 75 160.315 ;
      RECT 14.8 160.315 75 160.385 ;
      RECT 14.87 160.385 75 160.455 ;
      RECT 14.94 160.455 75 160.525 ;
      RECT 15.01 160.525 75 160.595 ;
      RECT 15.08 160.595 75 160.665 ;
      RECT 15.125 160.665 75 160.71 ;
      RECT 15.125 153.91 75 153.98 ;
      RECT 15.055 153.98 75 154.05 ;
      RECT 14.985 154.05 75 154.12 ;
      RECT 14.915 154.12 75 154.19 ;
      RECT 14.845 154.19 75 154.26 ;
      RECT 14.775 154.26 75 154.33 ;
      RECT 14.705 154.33 75 154.4 ;
      RECT 14.635 154.4 75 154.47 ;
      RECT 14.565 154.47 75 154.54 ;
      RECT 14.495 154.54 75 154.61 ;
      RECT 14.425 154.61 75 154.68 ;
      RECT 14.355 154.68 75 154.75 ;
      RECT 14.285 154.75 75 154.795 ;
      RECT 14.31 149.825 75 149.895 ;
      RECT 14.38 149.895 75 149.965 ;
      RECT 14.45 149.965 75 150.035 ;
      RECT 14.52 150.035 75 150.105 ;
      RECT 14.59 150.105 75 150.175 ;
      RECT 14.66 150.175 75 150.245 ;
      RECT 14.73 150.245 75 150.315 ;
      RECT 14.8 150.315 75 150.385 ;
      RECT 14.87 150.385 75 150.455 ;
      RECT 14.94 150.455 75 150.525 ;
      RECT 15.01 150.525 75 150.595 ;
      RECT 15.08 150.595 75 150.665 ;
      RECT 15.125 150.665 75 150.71 ;
      RECT 15.125 143.91 75 143.98 ;
      RECT 15.055 143.98 75 144.05 ;
      RECT 14.985 144.05 75 144.12 ;
      RECT 0 0 0.22 193.91 ;
      RECT 14.03 50.73 15.855 53.93 ;
      RECT 14.03 60.71 15.855 63.91 ;
      RECT 14.03 30.73 15.855 33.93 ;
      RECT 14.03 40.71 15.855 43.91 ;
      RECT 14.03 70.71 15.855 73.91 ;
      RECT 17.14 4.325 17.35 8.35 ;
      RECT 0 193.91 75 198 ;
      RECT 68.29 190.71 75 193.91 ;
      RECT 14.24 184.795 75 189.825 ;
      RECT 68.29 180.71 75 183.91 ;
      RECT 14.24 174.795 75 179.825 ;
      RECT 68.29 170.71 75 173.91 ;
      RECT 14.24 164.795 75 169.825 ;
      RECT 68.29 160.71 75 163.91 ;
      RECT 14.24 154.795 75 159.825 ;
      RECT 68.29 150.71 75 153.91 ;
      RECT 14.24 144.795 75 149.825 ;
      RECT 68.29 140.71 75 143.91 ;
      RECT 14.24 134.795 75 139.825 ;
      RECT 68.29 130.71 75 133.91 ;
      RECT 14.24 124.795 75 129.825 ;
      RECT 15.78 75.93 65.72 98.84 ;
      RECT 15.78 74.545 65.72 75.93 ;
      RECT 15.78 98.84 75 123.255 ;
      RECT 68.29 74.545 75 98.84 ;
      RECT 14.03 64.795 65.715 69.825 ;
      RECT 14.03 54.8 65.715 59.825 ;
      RECT 14.03 44.785 65.72 49.84 ;
      RECT 14.03 34.805 65.72 39.82 ;
      RECT 14.03 25.555 65.72 29.765 ;
      RECT 10.705 7.05 11.735 7.055 ;
      RECT 10.705 8.595 11.735 8.6 ;
      RECT 10.71 8.6 11.735 8.605 ;
      RECT 10.93 6.825 11.51 6.895 ;
      RECT 10.86 6.895 11.58 6.965 ;
      RECT 10.79 6.965 11.65 7.035 ;
      RECT 10.72 7.035 11.72 7.05 ;
      RECT 10.78 8.605 11.665 8.675 ;
      RECT 10.85 8.675 11.595 8.745 ;
      RECT 10.92 8.745 11.525 8.815 ;
      RECT 10.93 8.815 11.515 8.825 ;
      RECT 14.1 74.18 65.35 74.25 ;
      RECT 14.17 74.25 65.425 74.32 ;
      RECT 14.24 74.32 65.495 74.39 ;
      RECT 14.31 74.39 65.565 74.46 ;
      RECT 14.38 74.46 65.635 74.53 ;
      RECT 14.395 74.53 65.705 74.545 ;
      RECT 14.03 73.91 65.085 73.98 ;
      RECT 14.03 73.98 65.155 74.05 ;
      RECT 14.03 74.05 65.225 74.12 ;
      RECT 14.03 74.12 65.295 74.18 ;
      RECT 14.465 74.545 65.72 74.615 ;
      RECT 14.535 74.615 65.72 74.685 ;
      RECT 14.605 74.685 65.72 74.755 ;
      RECT 14.675 74.755 65.72 74.825 ;
      RECT 14.745 74.825 65.72 74.895 ;
      RECT 14.815 74.895 65.72 74.965 ;
      RECT 14.885 74.965 65.72 75.035 ;
      RECT 14.955 75.035 65.72 75.105 ;
      RECT 15.025 75.105 65.72 75.175 ;
      RECT 15.095 75.175 65.72 75.245 ;
      RECT 15.165 75.245 65.72 75.315 ;
      RECT 15.235 75.315 65.72 75.385 ;
      RECT 15.305 75.385 65.72 75.455 ;
      RECT 15.375 75.455 65.72 75.525 ;
      RECT 15.445 75.525 65.72 75.595 ;
      RECT 15.515 75.595 65.72 75.665 ;
      RECT 15.585 75.665 65.72 75.735 ;
      RECT 15.655 75.735 65.72 75.805 ;
      RECT 15.725 75.805 65.72 75.875 ;
      RECT 15.78 75.875 65.72 75.93 ;
      RECT 17.21 8.35 17.35 8.42 ;
      RECT 17.28 8.42 17.35 8.49 ;
      RECT 17.28 4.185 17.35 4.255 ;
      RECT 17.21 4.255 17.35 4.325 ;
      RECT 20.775 0.69 21.42 0.76 ;
      RECT 20.705 0.76 21.35 0.83 ;
      RECT 20.635 0.83 21.28 0.9 ;
      RECT 20.565 0.9 21.21 0.97 ;
      RECT 20.495 0.97 21.14 1.04 ;
      RECT 20.425 1.04 21.07 1.11 ;
      RECT 20.355 1.11 21.0 1.18 ;
      RECT 20.285 1.18 20.93 1.25 ;
      RECT 20.215 1.25 20.86 1.32 ;
      RECT 20.145 1.32 20.82 1.36 ;
      RECT 20.775 0 22.11 0.07 ;
      RECT 20.775 0.07 22.04 0.14 ;
      RECT 20.775 0.14 21.97 0.21 ;
      RECT 20.775 0.21 21.9 0.28 ;
      RECT 20.775 0.28 21.83 0.35 ;
      RECT 20.775 0.35 21.76 0.42 ;
      RECT 20.775 0.42 21.69 0.49 ;
      RECT 20.775 0.49 21.62 0.56 ;
      RECT 20.775 0.56 21.55 0.63 ;
      RECT 20.775 0.63 21.49 0.69 ;
      RECT 53.815 7.07 53.885 7.14 ;
      RECT 53.815 7.14 53.955 7.21 ;
      RECT 53.815 7.21 54.025 7.28 ;
      RECT 53.815 7.28 54.095 7.35 ;
      RECT 53.815 7.35 54.165 7.42 ;
      RECT 53.815 7.42 54.235 7.49 ;
      RECT 53.815 7.49 54.305 7.56 ;
      RECT 53.815 7.56 54.375 7.63 ;
      RECT 53.815 7.63 54.445 7.7 ;
      RECT 53.815 7.7 54.515 7.77 ;
      RECT 53.815 7.77 54.585 7.84 ;
      RECT 53.815 7.84 54.655 7.91 ;
      RECT 53.815 7.91 54.725 7.98 ;
      RECT 53.815 7.98 54.795 8.05 ;
      RECT 53.815 8.05 54.865 8.12 ;
      RECT 53.815 8.12 54.935 8.19 ;
      RECT 53.815 8.19 55.005 8.26 ;
      RECT 53.815 8.26 55.075 8.33 ;
      RECT 53.815 8.33 55.145 8.4 ;
      RECT 53.815 8.4 55.215 8.47 ;
      RECT 53.815 8.47 55.285 8.54 ;
      RECT 53.815 8.54 55.355 8.61 ;
      RECT 53.815 8.61 55.425 8.68 ;
      RECT 53.815 8.68 55.495 8.75 ;
      RECT 10.7 7.055 11.735 8.595 ;
    LAYER met1 ;
      RECT 0 18.49 75 198 ;
      RECT 0 0 15.185 1.27 ;
      RECT 0 1.27 8.215 18.49 ;
      RECT 9.265 15.255 16.19 15.525 ;
      RECT 9.265 15.2 16.46 15.255 ;
      RECT 9.265 3.345 16.515 15.2 ;
      RECT 9.335 3.28 16.515 3.345 ;
      RECT 9.535 3.08 16.515 3.28 ;
      RECT 16.245 16.83 75 18.49 ;
      RECT 17.125 15.955 75 16.83 ;
      RECT 17.205 15.875 36.025 15.955 ;
      RECT 17.205 2.055 36.025 15.875 ;
      RECT 17.685 1.58 36.025 2.055 ;
      RECT 17.845 1.42 36.025 1.58 ;
      RECT 37.265 1.51 56.015 1.58 ;
      RECT 37.195 1.58 56.015 15.955 ;
      RECT 37.355 1.42 56.015 1.51 ;
      RECT 56.705 0 75 15.955 ;
      RECT 17.7 1.705 35.885 1.775 ;
      RECT 17.63 1.775 35.885 1.78 ;
      RECT 17.845 1.56 35.81 1.6 ;
      RECT 17.805 1.6 35.85 1.635 ;
      RECT 17.925 1.48 18.825 1.52 ;
      RECT 17.885 1.52 18.865 1.56 ;
      RECT 19.985 1.48 20.885 1.52 ;
      RECT 19.945 1.52 20.925 1.56 ;
      RECT 22.045 1.48 22.945 1.52 ;
      RECT 22.005 1.52 22.985 1.56 ;
      RECT 24.105 1.48 25.005 1.52 ;
      RECT 24.065 1.52 25.045 1.56 ;
      RECT 26.165 1.48 27.065 1.52 ;
      RECT 26.125 1.52 27.105 1.56 ;
      RECT 28.225 1.48 29.125 1.52 ;
      RECT 28.185 1.52 29.165 1.56 ;
      RECT 30.285 1.48 31.185 1.52 ;
      RECT 30.245 1.52 31.225 1.56 ;
      RECT 32.345 1.48 33.245 1.52 ;
      RECT 32.305 1.52 33.285 1.56 ;
      RECT 34.405 1.48 35.305 1.52 ;
      RECT 34.365 1.52 35.345 1.56 ;
      RECT 37.41 1.56 55.875 1.6 ;
      RECT 37.37 1.6 55.875 1.635 ;
      RECT 37.915 1.48 38.815 1.52 ;
      RECT 37.875 1.52 38.855 1.56 ;
      RECT 39.975 1.48 40.875 1.52 ;
      RECT 39.935 1.52 40.915 1.56 ;
      RECT 42.035 1.48 42.935 1.52 ;
      RECT 41.995 1.52 42.975 1.56 ;
      RECT 44.095 1.48 44.995 1.52 ;
      RECT 44.055 1.52 45.035 1.56 ;
      RECT 46.155 1.48 47.055 1.52 ;
      RECT 46.115 1.52 47.095 1.56 ;
      RECT 48.215 1.48 49.115 1.52 ;
      RECT 48.175 1.52 49.155 1.56 ;
      RECT 50.275 1.48 51.175 1.52 ;
      RECT 50.235 1.52 51.215 1.56 ;
      RECT 52.335 1.48 53.235 1.52 ;
      RECT 52.295 1.52 53.275 1.56 ;
      RECT 54.395 1.48 55.295 1.52 ;
      RECT 54.355 1.52 55.335 1.56 ;
      RECT 20.345 17.175 32.885 17.245 ;
      RECT 20.275 17.245 32.885 17.315 ;
      RECT 20.205 17.315 32.885 17.385 ;
      RECT 20.135 17.385 32.885 17.455 ;
      RECT 20.065 17.455 32.885 17.525 ;
      RECT 19.995 17.525 32.885 17.595 ;
      RECT 19.925 17.595 32.885 17.665 ;
      RECT 19.855 17.665 32.885 17.735 ;
      RECT 19.785 17.735 32.885 17.805 ;
      RECT 19.715 17.805 32.885 17.875 ;
      RECT 19.645 17.875 32.885 17.945 ;
      RECT 19.575 17.945 32.885 18.015 ;
      RECT 19.505 18.015 32.885 18.085 ;
      RECT 19.435 18.085 32.885 18.135 ;
      RECT 20.345 17.175 32.885 17.245 ;
      RECT 20.275 17.245 32.885 17.315 ;
      RECT 20.205 17.315 32.885 17.385 ;
      RECT 20.135 17.385 32.885 17.455 ;
      RECT 20.065 17.455 32.885 17.525 ;
      RECT 19.995 17.525 32.885 17.595 ;
      RECT 19.925 17.595 32.885 17.665 ;
      RECT 19.855 17.665 32.885 17.735 ;
      RECT 19.785 17.735 32.885 17.805 ;
      RECT 19.715 17.805 32.885 17.875 ;
      RECT 19.645 17.875 32.885 17.945 ;
      RECT 19.575 17.945 32.885 18.015 ;
      RECT 19.505 18.015 32.885 18.085 ;
      RECT 19.435 18.085 32.885 18.135 ;
      RECT 9.405 3.335 16.375 15.2 ;
      RECT 12.405 6.22 13.375 12.385 ;
      RECT 9.475 15.2 16.25 15.27 ;
      RECT 9.545 15.27 16.18 15.34 ;
      RECT 9.59 15.34 16.135 15.385 ;
      RECT 9.59 3.22 16.26 3.28 ;
      RECT 9.53 3.28 16.32 3.335 ;
      RECT 8.075 18.63 17.345 21.635 ;
      RECT 8.075 194.995 17.345 198 ;
      RECT 16.385 16.89 17.345 18.63 ;
      RECT 17.625 1.78 35.885 1.835 ;
      RECT 35.885 16.89 40.335 21.635 ;
      RECT 35.885 194.995 75 198 ;
      RECT 37.335 4.64 40.34 16.89 ;
      RECT 37.335 1.635 55.875 4.64 ;
      RECT 52.87 4.64 55.875 16.89 ;
      RECT 52.875 16.89 59.845 21.635 ;
      RECT 56.845 3.005 59.85 16.89 ;
      RECT 56.845 0 75 3.005 ;
      RECT 71.995 18.63 75 194.995 ;
      RECT 71.995 3.005 75 16.89 ;
      RECT 72.0 16.89 75 18.63 ;
      RECT 0 0 8.075 198 ;
      RECT 3.0 3.002 5.075 21.63 ;
      RECT 3.0 21.63 72.0 195.0 ;
      RECT 19.385 18.135 32.885 19.095 ;
      RECT 19.385 19.095 72.0 21.63 ;
      RECT 17.345 2.115 35.885 198 ;
      RECT 20.345 4.56 32.885 17.175 ;
      RECT 40.335 4.56 52.875 19.095 ;
      RECT 59.845 3.0 72.0 19.095 ;
      RECT 0 0 16.19 0.07 ;
      RECT 0 0.07 16.12 0.14 ;
      RECT 0 0.14 16.05 0.21 ;
      RECT 0 0.21 15.98 0.28 ;
      RECT 0 0.28 15.91 0.35 ;
      RECT 0 0.35 15.84 0.42 ;
      RECT 0 0.42 15.77 0.49 ;
      RECT 0 0.49 15.7 0.56 ;
      RECT 0 0.56 15.63 0.63 ;
      RECT 0 0.63 15.56 0.7 ;
      RECT 0 0.7 15.49 0.77 ;
      RECT 0 0.77 15.42 0.84 ;
      RECT 0 0.84 15.35 0.91 ;
      RECT 0 0.91 15.28 0.98 ;
      RECT 0 0.98 15.21 1.05 ;
      RECT 0 1.05 15.14 1.12 ;
      RECT 0 1.12 15.13 1.13 ;
      RECT 17.18 16.095 75 16.165 ;
      RECT 17.11 16.165 75 16.235 ;
      RECT 17.04 16.235 75 16.305 ;
      RECT 16.97 16.305 75 16.375 ;
      RECT 16.9 16.375 75 16.445 ;
      RECT 16.83 16.445 75 16.515 ;
      RECT 16.76 16.515 75 16.585 ;
      RECT 16.69 16.585 75 16.655 ;
      RECT 16.62 16.655 75 16.725 ;
      RECT 16.55 16.725 75 16.795 ;
      RECT 16.48 16.795 75 16.865 ;
      RECT 16.41 16.865 75 16.89 ;
      RECT 17.345 15.93 35.885 16 ;
      RECT 17.275 16 35.885 16.07 ;
      RECT 17.205 16.07 35.885 16.095 ;
      RECT 17.625 1.835 35.885 1.905 ;
      RECT 17.555 1.905 35.885 1.975 ;
      RECT 17.485 1.975 35.885 2.045 ;
      RECT 17.415 2.045 35.885 2.115 ;
      RECT 17.77 1.635 35.885 1.705 ;
    LAYER li1 ;
      RECT 53.56 186.9 54.09 193.57 ;
      RECT 53.57 193.57 54.08 193.63 ;
      RECT 53.57 186.84 54.08 186.9 ;
      RECT 53.56 176.9 54.09 183.57 ;
      RECT 53.57 183.57 54.08 183.63 ;
      RECT 53.57 176.84 54.08 176.9 ;
      RECT 57.535 176.84 58.425 183.63 ;
      RECT 57.535 186.84 58.425 193.63 ;
      RECT 56.33 186.9 56.86 193.57 ;
      RECT 56.34 193.57 56.85 193.63 ;
      RECT 56.34 186.84 56.85 186.9 ;
      RECT 59.1 186.9 59.63 193.57 ;
      RECT 59.11 193.57 59.62 193.63 ;
      RECT 59.11 186.84 59.62 186.9 ;
      RECT 59.1 176.9 59.63 183.57 ;
      RECT 59.11 183.57 59.62 183.63 ;
      RECT 59.11 176.84 59.62 176.9 ;
      RECT 56.33 176.9 56.86 183.57 ;
      RECT 56.34 183.57 56.85 183.63 ;
      RECT 56.34 176.84 56.85 176.9 ;
      RECT 63.075 176.84 63.965 183.63 ;
      RECT 60.305 176.84 61.195 183.63 ;
      RECT 63.075 186.84 63.965 193.63 ;
      RECT 60.305 186.84 61.195 193.63 ;
      RECT 61.87 186.9 62.4 193.57 ;
      RECT 61.88 193.57 62.39 193.63 ;
      RECT 61.88 186.84 62.39 186.9 ;
      RECT 61.87 176.9 62.4 183.57 ;
      RECT 61.88 183.57 62.39 183.63 ;
      RECT 61.88 176.84 62.39 176.9 ;
      RECT 65.845 176.84 66.735 183.63 ;
      RECT 65.845 186.84 66.735 193.63 ;
      RECT 64.64 176.9 65.17 183.57 ;
      RECT 64.65 183.57 65.16 183.63 ;
      RECT 64.65 176.84 65.16 176.9 ;
      RECT 64.64 186.9 65.17 193.57 ;
      RECT 64.65 193.57 65.16 193.63 ;
      RECT 64.65 186.84 65.16 186.9 ;
      RECT 73.875 196.92 74.755 197.78 ;
      RECT 68.335 9.32 72.655 9.49 ;
      RECT 68.335 1.67 72.655 1.84 ;
      RECT 2.07 1.61 6.39 1.78 ;
      RECT 2.07 9.26 6.39 9.43 ;
      RECT 12.975 81.045 66.655 81.215 ;
      RECT 24.67 117.14 66.655 117.31 ;
      RECT 24.615 98.54 66.655 98.71 ;
      RECT 24.67 118.315 66.655 118.485 ;
      RECT 24.615 90.045 66.655 90.215 ;
      RECT 24.67 108.645 66.655 108.815 ;
      RECT 14.36 194.1 65.59 194.27 ;
      RECT 59.755 156.9 60.285 163.57 ;
      RECT 59.765 163.57 60.275 163.63 ;
      RECT 59.765 156.84 60.275 156.9 ;
      RECT 65.845 166.84 66.735 173.63 ;
      RECT 65.845 156.84 66.735 163.63 ;
      RECT 63.935 166.9 64.465 173.57 ;
      RECT 63.945 173.57 64.455 173.63 ;
      RECT 63.945 166.84 64.455 166.9 ;
      RECT 63.935 156.9 64.465 163.57 ;
      RECT 63.945 163.57 64.455 163.63 ;
      RECT 63.945 156.84 64.455 156.9 ;
      RECT 8.34 195.85 8.67 196.42 ;
      RECT 13.215 186.84 14.105 193.63 ;
      RECT 12.43 184.1 66.575 184.14 ;
      RECT 12.405 184.14 66.575 186.62 ;
      RECT 13.335 174.1 65.59 176.62 ;
      RECT 15.985 176.84 16.875 183.63 ;
      RECT 15.985 186.84 16.875 193.63 ;
      RECT 14.78 186.9 15.31 193.57 ;
      RECT 14.79 193.57 15.3 193.63 ;
      RECT 14.79 186.84 15.3 186.9 ;
      RECT 18.755 176.84 19.645 183.63 ;
      RECT 18.755 186.84 19.645 193.63 ;
      RECT 20.32 186.9 20.85 193.57 ;
      RECT 20.33 193.57 20.84 193.63 ;
      RECT 20.33 186.84 20.84 186.9 ;
      RECT 17.55 186.9 18.08 193.57 ;
      RECT 17.56 193.57 18.07 193.63 ;
      RECT 17.56 186.84 18.07 186.9 ;
      RECT 20.32 176.9 20.85 183.57 ;
      RECT 20.33 183.57 20.84 183.63 ;
      RECT 20.33 176.84 20.84 176.9 ;
      RECT 17.55 176.9 18.08 183.57 ;
      RECT 17.56 183.57 18.07 183.63 ;
      RECT 17.56 176.84 18.07 176.9 ;
      RECT 24.295 176.84 25.185 183.63 ;
      RECT 21.525 176.84 22.415 183.63 ;
      RECT 24.295 186.84 25.185 193.63 ;
      RECT 21.525 186.84 22.415 193.63 ;
      RECT 23.09 176.9 23.62 183.57 ;
      RECT 23.1 183.57 23.61 183.63 ;
      RECT 23.1 176.84 23.61 176.9 ;
      RECT 23.09 186.9 23.62 193.57 ;
      RECT 23.1 193.57 23.61 193.63 ;
      RECT 23.1 186.84 23.61 186.9 ;
      RECT 27.065 176.84 27.955 183.63 ;
      RECT 27.065 186.84 27.955 193.63 ;
      RECT 28.63 176.9 29.16 183.57 ;
      RECT 28.64 183.57 29.15 183.63 ;
      RECT 28.64 176.84 29.15 176.9 ;
      RECT 25.86 176.9 26.39 183.57 ;
      RECT 25.87 183.57 26.38 183.63 ;
      RECT 25.87 176.84 26.38 176.9 ;
      RECT 28.63 186.9 29.16 193.57 ;
      RECT 28.64 193.57 29.15 193.63 ;
      RECT 28.64 186.84 29.15 186.9 ;
      RECT 25.86 186.9 26.39 193.57 ;
      RECT 25.87 193.57 26.38 193.63 ;
      RECT 25.87 186.84 26.38 186.9 ;
      RECT 29.835 176.84 30.725 183.63 ;
      RECT 29.835 186.84 30.725 193.63 ;
      RECT 31.4 176.9 31.93 183.57 ;
      RECT 31.41 183.57 31.92 183.63 ;
      RECT 31.41 176.84 31.92 176.9 ;
      RECT 31.4 186.9 31.93 193.57 ;
      RECT 31.41 193.57 31.92 193.63 ;
      RECT 31.41 186.84 31.92 186.9 ;
      RECT 35.375 176.84 36.265 183.63 ;
      RECT 32.605 176.84 33.495 183.63 ;
      RECT 35.375 186.84 36.265 193.63 ;
      RECT 32.605 186.84 33.495 193.63 ;
      RECT 34.17 186.9 34.7 193.57 ;
      RECT 34.18 193.57 34.69 193.63 ;
      RECT 34.18 186.84 34.69 186.9 ;
      RECT 34.17 176.9 34.7 183.57 ;
      RECT 34.18 183.57 34.69 183.63 ;
      RECT 34.18 176.84 34.69 176.9 ;
      RECT 38.145 176.84 39.035 183.63 ;
      RECT 38.145 186.84 39.035 193.63 ;
      RECT 36.94 176.9 37.47 183.57 ;
      RECT 36.95 183.57 37.46 183.63 ;
      RECT 36.95 176.84 37.46 176.9 ;
      RECT 36.94 186.9 37.47 193.57 ;
      RECT 36.95 193.57 37.46 193.63 ;
      RECT 36.95 186.84 37.46 186.9 ;
      RECT 39.71 176.9 40.24 183.57 ;
      RECT 39.72 183.57 40.23 183.63 ;
      RECT 39.72 176.84 40.23 176.9 ;
      RECT 39.71 186.9 40.24 193.57 ;
      RECT 39.72 193.57 40.23 193.63 ;
      RECT 39.72 186.84 40.23 186.9 ;
      RECT 43.685 176.84 44.575 183.63 ;
      RECT 40.915 176.84 41.805 183.63 ;
      RECT 43.685 186.84 44.575 193.63 ;
      RECT 40.915 186.84 41.805 193.63 ;
      RECT 42.48 176.9 43.01 183.57 ;
      RECT 42.49 183.57 43 183.63 ;
      RECT 42.49 176.84 43 176.9 ;
      RECT 42.48 186.9 43.01 193.57 ;
      RECT 42.49 193.57 43 193.63 ;
      RECT 42.49 186.84 43 186.9 ;
      RECT 46.455 176.84 47.345 183.63 ;
      RECT 46.455 186.84 47.345 193.63 ;
      RECT 45.25 176.9 45.78 183.57 ;
      RECT 45.26 183.57 45.77 183.63 ;
      RECT 45.26 176.84 45.77 176.9 ;
      RECT 45.25 186.9 45.78 193.57 ;
      RECT 45.26 193.57 45.77 193.63 ;
      RECT 45.26 186.84 45.77 186.9 ;
      RECT 49.225 176.84 50.115 183.63 ;
      RECT 49.225 186.84 50.115 193.63 ;
      RECT 48.02 176.9 48.55 183.57 ;
      RECT 48.03 183.57 48.54 183.63 ;
      RECT 48.03 176.84 48.54 176.9 ;
      RECT 50.79 176.9 51.32 183.57 ;
      RECT 50.8 183.57 51.31 183.63 ;
      RECT 50.8 176.84 51.31 176.9 ;
      RECT 50.79 186.9 51.32 193.57 ;
      RECT 50.8 193.57 51.31 193.63 ;
      RECT 50.8 186.84 51.31 186.9 ;
      RECT 48.02 186.9 48.55 193.57 ;
      RECT 48.03 193.57 48.54 193.63 ;
      RECT 48.03 186.84 48.54 186.9 ;
      RECT 54.765 176.84 55.655 183.63 ;
      RECT 51.995 176.84 52.885 183.63 ;
      RECT 54.765 186.84 55.655 193.63 ;
      RECT 51.995 186.84 52.885 193.63 ;
      RECT 53.305 136.84 54.195 143.63 ;
      RECT 53.305 146.84 54.195 153.63 ;
      RECT 55.575 136.9 56.105 143.57 ;
      RECT 55.585 143.57 56.095 143.63 ;
      RECT 55.585 136.84 56.095 136.9 ;
      RECT 55.575 146.9 56.105 153.57 ;
      RECT 55.585 153.57 56.095 153.63 ;
      RECT 55.585 146.84 56.095 146.9 ;
      RECT 55.575 128.73 56.105 133.925 ;
      RECT 57.485 128.735 58.375 133.485 ;
      RECT 57.665 133.485 58.195 133.755 ;
      RECT 57.665 128.73 58.195 128.735 ;
      RECT 57.485 136.84 58.375 143.63 ;
      RECT 57.485 146.84 58.375 153.63 ;
      RECT 61.665 128.735 62.555 133.485 ;
      RECT 61.845 133.485 62.375 133.755 ;
      RECT 61.845 128.73 62.375 128.735 ;
      RECT 61.665 136.84 62.555 143.63 ;
      RECT 61.665 146.84 62.555 153.63 ;
      RECT 59.755 136.9 60.285 143.57 ;
      RECT 59.765 143.57 60.275 143.63 ;
      RECT 59.765 136.84 60.275 136.9 ;
      RECT 59.755 146.9 60.285 153.57 ;
      RECT 59.765 153.57 60.275 153.63 ;
      RECT 59.765 146.84 60.275 146.9 ;
      RECT 59.755 128.73 60.285 133.925 ;
      RECT 65.845 128.735 66.735 133.485 ;
      RECT 66.025 133.485 66.555 133.755 ;
      RECT 66.025 128.73 66.555 128.735 ;
      RECT 65.845 136.84 66.735 143.63 ;
      RECT 65.845 146.84 66.735 153.63 ;
      RECT 63.935 136.9 64.465 143.57 ;
      RECT 63.945 143.57 64.455 143.63 ;
      RECT 63.945 136.84 64.455 136.9 ;
      RECT 63.935 146.9 64.465 153.57 ;
      RECT 63.945 153.57 64.455 153.63 ;
      RECT 63.945 146.84 64.455 146.9 ;
      RECT 63.935 128.73 64.465 133.925 ;
      RECT 13.365 154.1 65.59 156.62 ;
      RECT 13.365 164.1 65.59 166.62 ;
      RECT 15.685 156.84 16.575 163.63 ;
      RECT 15.685 166.84 16.575 173.63 ;
      RECT 19.865 156.84 20.755 163.63 ;
      RECT 19.865 166.84 20.755 173.63 ;
      RECT 17.955 166.9 18.485 173.57 ;
      RECT 17.965 173.57 18.475 173.63 ;
      RECT 17.965 166.84 18.475 166.9 ;
      RECT 17.955 156.9 18.485 163.57 ;
      RECT 17.965 163.57 18.475 163.63 ;
      RECT 17.965 156.84 18.475 156.9 ;
      RECT 24.045 156.84 24.935 163.63 ;
      RECT 24.045 166.84 24.935 173.63 ;
      RECT 22.135 166.9 22.665 173.57 ;
      RECT 22.145 173.57 22.655 173.63 ;
      RECT 22.145 166.84 22.655 166.9 ;
      RECT 22.135 156.9 22.665 163.57 ;
      RECT 22.145 163.57 22.655 163.63 ;
      RECT 22.145 156.84 22.655 156.9 ;
      RECT 28.225 156.84 29.115 163.63 ;
      RECT 28.225 166.84 29.115 173.63 ;
      RECT 26.315 166.9 26.845 173.57 ;
      RECT 26.325 173.57 26.835 173.63 ;
      RECT 26.325 166.84 26.835 166.9 ;
      RECT 26.315 156.9 26.845 163.57 ;
      RECT 26.325 163.57 26.835 163.63 ;
      RECT 26.325 156.84 26.835 156.9 ;
      RECT 32.405 156.84 33.295 163.63 ;
      RECT 32.405 166.84 33.295 173.63 ;
      RECT 30.495 166.9 31.025 173.57 ;
      RECT 30.505 173.57 31.015 173.63 ;
      RECT 30.505 166.84 31.015 166.9 ;
      RECT 30.495 156.9 31.025 163.57 ;
      RECT 30.505 163.57 31.015 163.63 ;
      RECT 30.505 156.84 31.015 156.9 ;
      RECT 34.675 166.9 35.205 173.57 ;
      RECT 34.685 173.57 35.195 173.63 ;
      RECT 34.685 166.84 35.195 166.9 ;
      RECT 34.675 156.9 35.205 163.57 ;
      RECT 34.685 163.57 35.195 163.63 ;
      RECT 34.685 156.84 35.195 156.9 ;
      RECT 36.585 156.84 37.475 163.63 ;
      RECT 36.585 166.84 37.475 173.63 ;
      RECT 38.855 166.9 39.385 173.57 ;
      RECT 38.865 173.57 39.375 173.63 ;
      RECT 38.865 166.84 39.375 166.9 ;
      RECT 38.855 156.9 39.385 163.57 ;
      RECT 38.865 163.57 39.375 163.63 ;
      RECT 38.865 156.84 39.375 156.9 ;
      RECT 40.765 156.84 41.655 163.63 ;
      RECT 40.765 166.84 41.655 173.63 ;
      RECT 43.035 166.9 43.565 173.57 ;
      RECT 43.045 173.57 43.555 173.63 ;
      RECT 43.045 166.84 43.555 166.9 ;
      RECT 43.035 156.9 43.565 163.57 ;
      RECT 43.045 163.57 43.555 163.63 ;
      RECT 43.045 156.84 43.555 156.9 ;
      RECT 44.945 156.84 45.835 163.63 ;
      RECT 44.945 166.84 45.835 173.63 ;
      RECT 47.215 166.9 47.745 173.57 ;
      RECT 47.225 173.57 47.735 173.63 ;
      RECT 47.225 166.84 47.735 166.9 ;
      RECT 47.215 156.9 47.745 163.57 ;
      RECT 47.225 163.57 47.735 163.63 ;
      RECT 47.225 156.84 47.735 156.9 ;
      RECT 49.125 156.84 50.015 163.63 ;
      RECT 49.125 166.84 50.015 173.63 ;
      RECT 51.395 166.9 51.925 173.57 ;
      RECT 51.405 173.57 51.915 173.63 ;
      RECT 51.405 166.84 51.915 166.9 ;
      RECT 51.395 156.9 51.925 163.57 ;
      RECT 51.405 163.57 51.915 163.63 ;
      RECT 51.405 156.84 51.915 156.9 ;
      RECT 53.305 156.84 54.195 163.63 ;
      RECT 53.305 166.84 54.195 173.63 ;
      RECT 55.575 166.9 56.105 173.57 ;
      RECT 55.585 173.57 56.095 173.63 ;
      RECT 55.585 166.84 56.095 166.9 ;
      RECT 55.575 156.9 56.105 163.57 ;
      RECT 55.585 163.57 56.095 163.63 ;
      RECT 55.585 156.84 56.095 156.9 ;
      RECT 57.485 156.84 58.375 163.63 ;
      RECT 57.485 166.84 58.375 173.63 ;
      RECT 61.665 166.84 62.555 173.63 ;
      RECT 61.665 156.84 62.555 163.63 ;
      RECT 59.755 166.9 60.285 173.57 ;
      RECT 59.765 173.57 60.275 173.63 ;
      RECT 59.765 166.84 60.275 166.9 ;
      RECT 23.805 115.55 24.215 116.67 ;
      RECT 23.635 109.88 24.215 115.55 ;
      RECT 23.635 101.385 24.215 108.175 ;
      RECT 25.31 110.45 25.535 115.33 ;
      RECT 25.31 115.33 25.48 116.67 ;
      RECT 25.31 109.88 25.48 110.45 ;
      RECT 25.31 120.08 25.535 124.86 ;
      RECT 25.31 124.86 25.48 125.745 ;
      RECT 25.31 118.955 25.48 120.08 ;
      RECT 25.31 101.385 25.535 106.255 ;
      RECT 25.31 106.255 25.48 108.175 ;
      RECT 33.59 109.88 33.76 116.67 ;
      RECT 33.59 120.08 33.765 124.86 ;
      RECT 33.59 124.86 33.76 125.745 ;
      RECT 33.59 118.955 33.76 120.08 ;
      RECT 33.59 101.385 33.76 108.175 ;
      RECT 41.87 109.88 42.04 116.67 ;
      RECT 41.87 118.955 42.04 125.745 ;
      RECT 41.87 101.385 42.04 108.175 ;
      RECT 50.15 109.88 50.32 116.67 ;
      RECT 50.15 118.955 50.32 125.745 ;
      RECT 50.15 101.385 50.32 108.175 ;
      RECT 58.43 109.88 58.6 116.67 ;
      RECT 58.43 118.955 58.6 125.745 ;
      RECT 58.43 101.385 58.6 108.175 ;
      RECT 66.71 109.88 66.88 116.67 ;
      RECT 66.71 118.955 66.88 125.745 ;
      RECT 66.71 101.385 66.88 108.175 ;
      RECT 13.365 145.62 65.59 146.62 ;
      RECT 23.405 144.1 65.59 145.62 ;
      RECT 13.365 145.615 14.305 145.62 ;
      RECT 15.685 146.84 16.575 153.63 ;
      RECT 19.865 146.84 20.755 153.63 ;
      RECT 17.955 146.9 18.485 153.57 ;
      RECT 17.965 153.57 18.475 153.63 ;
      RECT 17.965 146.84 18.475 146.9 ;
      RECT 24.045 128.735 24.935 133.485 ;
      RECT 24.225 133.485 24.755 133.76 ;
      RECT 24.225 128.73 24.755 128.735 ;
      RECT 24.045 136.84 24.935 143.63 ;
      RECT 24.045 146.84 24.935 153.63 ;
      RECT 22.135 146.9 22.665 153.57 ;
      RECT 22.145 153.57 22.655 153.63 ;
      RECT 22.145 146.84 22.655 146.9 ;
      RECT 21.69 134.1 65.59 136.62 ;
      RECT 21.66 128.01 65.59 128.515 ;
      RECT 28.225 128.735 29.115 133.485 ;
      RECT 28.405 133.485 28.935 133.76 ;
      RECT 28.225 136.84 29.115 143.63 ;
      RECT 28.225 146.84 29.115 153.63 ;
      RECT 26.315 146.9 26.845 153.57 ;
      RECT 26.325 153.57 26.835 153.63 ;
      RECT 26.325 146.84 26.835 146.9 ;
      RECT 26.315 136.9 26.845 143.57 ;
      RECT 26.325 143.57 26.835 143.63 ;
      RECT 26.325 136.84 26.835 136.9 ;
      RECT 26.315 128.73 26.845 133.715 ;
      RECT 32.405 128.735 33.295 133.485 ;
      RECT 32.585 133.485 33.115 133.755 ;
      RECT 32.585 128.73 33.115 128.735 ;
      RECT 32.405 136.84 33.295 143.63 ;
      RECT 32.405 146.84 33.295 153.63 ;
      RECT 30.495 146.9 31.025 153.57 ;
      RECT 30.505 153.57 31.015 153.63 ;
      RECT 30.505 146.84 31.015 146.9 ;
      RECT 30.495 136.9 31.025 143.57 ;
      RECT 30.505 143.57 31.015 143.63 ;
      RECT 30.505 136.84 31.015 136.9 ;
      RECT 30.495 128.73 31.025 133.715 ;
      RECT 34.675 146.9 35.205 153.57 ;
      RECT 34.685 153.57 35.195 153.63 ;
      RECT 34.685 146.84 35.195 146.9 ;
      RECT 34.675 136.9 35.205 143.57 ;
      RECT 34.685 143.57 35.195 143.63 ;
      RECT 34.685 136.84 35.195 136.9 ;
      RECT 34.675 128.73 35.205 133.84 ;
      RECT 36.585 128.735 37.475 133.485 ;
      RECT 36.765 133.485 37.295 133.755 ;
      RECT 36.765 128.73 37.295 128.735 ;
      RECT 36.585 136.84 37.475 143.63 ;
      RECT 36.585 146.84 37.475 153.63 ;
      RECT 38.855 146.9 39.385 153.57 ;
      RECT 38.865 153.57 39.375 153.63 ;
      RECT 38.865 146.84 39.375 146.9 ;
      RECT 38.855 136.9 39.385 143.57 ;
      RECT 38.865 143.57 39.375 143.63 ;
      RECT 38.865 136.84 39.375 136.9 ;
      RECT 38.855 128.73 39.385 133.925 ;
      RECT 40.765 128.735 41.655 133.485 ;
      RECT 40.945 133.485 41.475 133.755 ;
      RECT 40.945 128.73 41.475 128.735 ;
      RECT 40.765 136.84 41.655 143.63 ;
      RECT 40.765 146.84 41.655 153.63 ;
      RECT 43.035 146.9 43.565 153.57 ;
      RECT 43.045 153.57 43.555 153.63 ;
      RECT 43.045 146.84 43.555 146.9 ;
      RECT 43.035 136.9 43.565 143.57 ;
      RECT 43.045 143.57 43.555 143.63 ;
      RECT 43.045 136.84 43.555 136.9 ;
      RECT 43.035 128.73 43.565 133.925 ;
      RECT 44.945 128.735 45.835 133.485 ;
      RECT 45.125 133.485 45.655 133.755 ;
      RECT 45.125 128.73 45.655 128.735 ;
      RECT 44.945 136.84 45.835 143.63 ;
      RECT 44.945 146.84 45.835 153.63 ;
      RECT 47.215 146.9 47.745 153.57 ;
      RECT 47.225 153.57 47.735 153.63 ;
      RECT 47.225 146.84 47.735 146.9 ;
      RECT 47.215 136.9 47.745 143.57 ;
      RECT 47.225 143.57 47.735 143.63 ;
      RECT 47.225 136.84 47.735 136.9 ;
      RECT 47.215 128.73 47.745 133.925 ;
      RECT 49.125 128.735 50.015 133.485 ;
      RECT 49.305 133.485 49.835 133.755 ;
      RECT 49.305 128.73 49.835 128.735 ;
      RECT 49.125 136.84 50.015 143.63 ;
      RECT 49.125 146.84 50.015 153.63 ;
      RECT 51.395 136.9 51.925 143.57 ;
      RECT 51.405 143.57 51.915 143.63 ;
      RECT 51.405 136.84 51.915 136.9 ;
      RECT 51.395 146.9 51.925 153.57 ;
      RECT 51.405 153.57 51.915 153.63 ;
      RECT 51.405 146.84 51.915 146.9 ;
      RECT 51.395 128.73 51.925 133.925 ;
      RECT 53.305 128.735 54.195 133.485 ;
      RECT 53.485 133.485 54.015 133.755 ;
      RECT 53.485 128.73 54.015 128.735 ;
      RECT 35.555 71.59 36.085 71.725 ;
      RECT 32.605 66.84 33.495 71.59 ;
      RECT 32.785 71.59 33.315 71.725 ;
      RECT 35.375 56.84 36.265 63.63 ;
      RECT 32.605 56.84 33.495 63.63 ;
      RECT 34.17 56.9 34.7 63.57 ;
      RECT 34.18 63.57 34.69 63.63 ;
      RECT 34.18 56.84 34.69 56.9 ;
      RECT 34.17 66.9 34.7 71.725 ;
      RECT 34.18 66.84 34.69 66.9 ;
      RECT 38.145 66.84 39.035 71.59 ;
      RECT 38.325 71.59 38.855 71.725 ;
      RECT 38.145 56.84 39.035 63.63 ;
      RECT 39.71 56.9 40.24 63.57 ;
      RECT 39.72 63.57 40.23 63.63 ;
      RECT 39.72 56.84 40.23 56.9 ;
      RECT 36.94 56.9 37.47 63.57 ;
      RECT 36.95 63.57 37.46 63.63 ;
      RECT 36.95 56.84 37.46 56.9 ;
      RECT 39.71 66.9 40.24 71.725 ;
      RECT 39.72 66.84 40.23 66.9 ;
      RECT 36.94 66.9 37.47 71.725 ;
      RECT 36.95 66.84 37.46 66.9 ;
      RECT 43.685 66.84 44.575 71.59 ;
      RECT 43.865 71.59 44.395 71.725 ;
      RECT 40.915 66.84 41.805 71.59 ;
      RECT 41.095 71.59 41.625 71.725 ;
      RECT 43.685 56.84 44.575 63.63 ;
      RECT 40.915 56.84 41.805 63.63 ;
      RECT 42.48 56.9 43.01 63.57 ;
      RECT 42.49 63.57 43 63.63 ;
      RECT 42.49 56.84 43 56.9 ;
      RECT 42.48 66.9 43.01 71.725 ;
      RECT 42.49 66.84 43 66.9 ;
      RECT 46.455 66.84 47.345 71.59 ;
      RECT 46.635 71.59 47.165 71.725 ;
      RECT 46.455 56.84 47.345 63.63 ;
      RECT 45.25 56.9 45.78 63.57 ;
      RECT 45.26 63.57 45.77 63.63 ;
      RECT 45.26 56.84 45.77 56.9 ;
      RECT 45.25 66.9 45.78 71.725 ;
      RECT 45.26 66.84 45.77 66.9 ;
      RECT 49.225 66.84 50.115 71.59 ;
      RECT 49.405 71.59 49.935 71.725 ;
      RECT 49.225 56.84 50.115 63.63 ;
      RECT 48.02 56.9 48.55 63.57 ;
      RECT 48.03 63.57 48.54 63.63 ;
      RECT 48.03 56.84 48.54 56.9 ;
      RECT 50.79 56.9 51.32 63.57 ;
      RECT 50.8 63.57 51.31 63.63 ;
      RECT 50.8 56.84 51.31 56.9 ;
      RECT 50.79 66.9 51.32 71.725 ;
      RECT 50.8 66.84 51.31 66.9 ;
      RECT 48.02 66.9 48.55 71.725 ;
      RECT 48.03 66.84 48.54 66.9 ;
      RECT 54.765 66.84 55.655 71.59 ;
      RECT 54.945 71.59 55.475 71.725 ;
      RECT 51.995 66.84 52.885 71.59 ;
      RECT 52.175 71.59 52.705 71.725 ;
      RECT 54.765 56.84 55.655 63.63 ;
      RECT 51.995 56.84 52.885 63.63 ;
      RECT 53.56 56.9 54.09 63.57 ;
      RECT 53.57 63.57 54.08 63.63 ;
      RECT 53.57 56.84 54.08 56.9 ;
      RECT 53.56 66.9 54.09 71.725 ;
      RECT 53.57 66.84 54.08 66.9 ;
      RECT 57.535 66.84 58.425 71.59 ;
      RECT 57.715 71.59 58.245 71.725 ;
      RECT 57.535 56.84 58.425 63.63 ;
      RECT 56.33 56.9 56.86 63.57 ;
      RECT 56.34 63.57 56.85 63.63 ;
      RECT 56.34 56.84 56.85 56.9 ;
      RECT 59.1 56.9 59.63 63.57 ;
      RECT 59.11 63.57 59.62 63.63 ;
      RECT 59.11 56.84 59.62 56.9 ;
      RECT 56.33 66.9 56.86 71.725 ;
      RECT 56.34 66.84 56.85 66.9 ;
      RECT 59.1 66.9 59.63 71.725 ;
      RECT 59.11 66.84 59.62 66.9 ;
      RECT 63.075 66.84 63.965 71.59 ;
      RECT 63.255 71.59 63.785 71.725 ;
      RECT 60.305 66.84 61.195 71.59 ;
      RECT 60.485 71.59 61.015 71.725 ;
      RECT 63.075 56.84 63.965 63.63 ;
      RECT 60.305 56.84 61.195 63.63 ;
      RECT 61.87 56.9 62.4 63.57 ;
      RECT 61.88 63.57 62.39 63.63 ;
      RECT 61.88 56.84 62.39 56.9 ;
      RECT 61.87 66.9 62.4 71.725 ;
      RECT 61.88 66.84 62.39 66.9 ;
      RECT 65.845 66.84 66.735 71.59 ;
      RECT 66.025 71.59 66.555 71.725 ;
      RECT 65.845 56.84 66.735 63.63 ;
      RECT 64.64 56.9 65.17 63.57 ;
      RECT 64.65 63.57 65.16 63.63 ;
      RECT 64.65 56.84 65.16 56.9 ;
      RECT 64.64 66.9 65.17 71.725 ;
      RECT 64.65 66.84 65.16 66.9 ;
      RECT 10.92 84.33 11.83 84.585 ;
      RECT 10.915 84.16 11.83 84.33 ;
      RECT 10.92 83.82 11.83 84.16 ;
      RECT 12.75 75.785 12.92 80.535 ;
      RECT 17.03 75.785 17.2 80.535 ;
      RECT 19.495 83.82 20.405 84.585 ;
      RECT 23.685 82.785 24.215 89.575 ;
      RECT 23.685 91.28 24.215 98.07 ;
      RECT 25.31 91.28 25.48 98.07 ;
      RECT 25.31 82.785 25.48 89.575 ;
      RECT 25.31 75.785 25.48 80.535 ;
      RECT 33.59 75.785 33.76 80.535 ;
      RECT 33.59 91.28 33.76 98.07 ;
      RECT 33.59 82.785 33.76 89.575 ;
      RECT 41.87 75.785 42.04 80.535 ;
      RECT 41.87 91.28 42.04 98.07 ;
      RECT 41.87 82.785 42.04 89.575 ;
      RECT 50.15 75.785 50.32 80.535 ;
      RECT 50.15 91.28 50.32 98.07 ;
      RECT 50.15 82.785 50.32 89.575 ;
      RECT 58.43 75.785 58.6 80.535 ;
      RECT 58.43 91.28 58.6 98.07 ;
      RECT 58.43 82.785 58.6 89.575 ;
      RECT 66.71 91.28 66.88 98.07 ;
      RECT 66.71 82.785 66.88 89.575 ;
      RECT 66.71 75.785 66.88 80.535 ;
      RECT 23.805 125.295 24.215 125.745 ;
      RECT 23.635 120.08 24.215 125.295 ;
      RECT 23.805 118.955 24.215 120.08 ;
      RECT 48.03 43.57 48.54 43.63 ;
      RECT 48.03 36.84 48.54 36.9 ;
      RECT 50.79 36.9 51.32 43.57 ;
      RECT 50.8 43.57 51.31 43.63 ;
      RECT 50.8 36.84 51.31 36.9 ;
      RECT 54.765 36.84 55.655 43.63 ;
      RECT 51.995 36.84 52.885 43.63 ;
      RECT 54.765 26.84 55.655 33.63 ;
      RECT 51.995 26.84 52.885 33.63 ;
      RECT 54.765 46.84 55.655 53.63 ;
      RECT 51.995 46.84 52.885 53.63 ;
      RECT 53.56 26.9 54.09 33.57 ;
      RECT 53.57 33.57 54.08 33.63 ;
      RECT 53.57 26.84 54.08 26.9 ;
      RECT 53.56 46.9 54.09 53.57 ;
      RECT 53.57 53.57 54.08 53.63 ;
      RECT 53.57 46.84 54.08 46.9 ;
      RECT 53.56 36.9 54.09 43.57 ;
      RECT 53.57 43.57 54.08 43.63 ;
      RECT 53.57 36.84 54.08 36.9 ;
      RECT 57.535 36.84 58.425 43.63 ;
      RECT 57.535 26.84 58.425 33.63 ;
      RECT 57.535 46.84 58.425 53.63 ;
      RECT 56.33 26.9 56.86 33.57 ;
      RECT 56.34 33.57 56.85 33.63 ;
      RECT 56.34 26.84 56.85 26.9 ;
      RECT 59.1 26.9 59.63 33.57 ;
      RECT 59.11 33.57 59.62 33.63 ;
      RECT 59.11 26.84 59.62 26.9 ;
      RECT 56.33 46.9 56.86 53.57 ;
      RECT 56.34 53.57 56.85 53.63 ;
      RECT 56.34 46.84 56.85 46.9 ;
      RECT 59.1 46.9 59.63 53.57 ;
      RECT 59.11 53.57 59.62 53.63 ;
      RECT 59.11 46.84 59.62 46.9 ;
      RECT 56.33 36.9 56.86 43.57 ;
      RECT 56.34 43.57 56.85 43.63 ;
      RECT 56.34 36.84 56.85 36.9 ;
      RECT 59.1 36.9 59.63 43.57 ;
      RECT 59.11 43.57 59.62 43.63 ;
      RECT 59.11 36.84 59.62 36.9 ;
      RECT 63.075 36.84 63.965 43.63 ;
      RECT 60.305 36.84 61.195 43.63 ;
      RECT 63.075 26.84 63.965 33.63 ;
      RECT 60.305 26.84 61.195 33.63 ;
      RECT 63.075 46.84 63.965 53.63 ;
      RECT 60.305 46.84 61.195 53.63 ;
      RECT 61.87 26.9 62.4 33.57 ;
      RECT 61.88 33.57 62.39 33.63 ;
      RECT 61.88 26.84 62.39 26.9 ;
      RECT 61.87 46.9 62.4 53.57 ;
      RECT 61.88 53.57 62.39 53.63 ;
      RECT 61.88 46.84 62.39 46.9 ;
      RECT 61.87 36.9 62.4 43.57 ;
      RECT 61.88 43.57 62.39 43.63 ;
      RECT 61.88 36.84 62.39 36.9 ;
      RECT 65.845 36.84 66.735 43.63 ;
      RECT 65.845 26.84 66.735 33.63 ;
      RECT 65.845 46.84 66.735 53.63 ;
      RECT 64.64 46.9 65.17 53.57 ;
      RECT 64.65 53.57 65.16 53.63 ;
      RECT 64.65 46.84 65.16 46.9 ;
      RECT 64.64 36.9 65.17 43.57 ;
      RECT 64.65 43.57 65.16 43.63 ;
      RECT 64.65 36.84 65.16 36.9 ;
      RECT 64.64 26.9 65.17 33.57 ;
      RECT 64.65 33.57 65.16 33.63 ;
      RECT 64.65 26.84 65.16 26.9 ;
      RECT 13.215 66.84 14.105 71.59 ;
      RECT 13.395 71.59 13.925 71.725 ;
      RECT 13.215 56.84 14.105 63.63 ;
      RECT 13.19 54.1 65.59 56.62 ;
      RECT 13.06 64.1 65.59 66.62 ;
      RECT 15.985 66.84 16.875 71.59 ;
      RECT 16.165 71.59 16.695 71.725 ;
      RECT 15.985 56.84 16.875 63.63 ;
      RECT 14.78 56.9 15.31 63.57 ;
      RECT 14.79 63.57 15.3 63.63 ;
      RECT 14.79 56.84 15.3 56.9 ;
      RECT 14.78 66.9 15.31 71.725 ;
      RECT 14.79 66.84 15.3 66.9 ;
      RECT 18.755 66.84 19.645 71.59 ;
      RECT 18.935 71.59 19.465 71.725 ;
      RECT 18.755 56.84 19.645 63.63 ;
      RECT 20.32 56.9 20.85 63.57 ;
      RECT 20.33 63.57 20.84 63.63 ;
      RECT 20.33 56.84 20.84 56.9 ;
      RECT 17.55 56.9 18.08 63.57 ;
      RECT 17.56 63.57 18.07 63.63 ;
      RECT 17.56 56.84 18.07 56.9 ;
      RECT 20.32 66.9 20.85 71.725 ;
      RECT 20.33 66.84 20.84 66.9 ;
      RECT 17.55 66.9 18.08 71.725 ;
      RECT 17.56 66.84 18.07 66.9 ;
      RECT 24.295 66.84 25.185 71.59 ;
      RECT 24.475 71.59 25.005 71.725 ;
      RECT 21.525 66.84 22.415 71.59 ;
      RECT 21.705 71.59 22.235 71.725 ;
      RECT 24.295 56.84 25.185 63.63 ;
      RECT 21.525 56.84 22.415 63.63 ;
      RECT 23.09 56.9 23.62 63.57 ;
      RECT 23.1 63.57 23.61 63.63 ;
      RECT 23.1 56.84 23.61 56.9 ;
      RECT 23.09 66.9 23.62 71.725 ;
      RECT 23.1 66.84 23.61 66.9 ;
      RECT 27.065 66.84 27.955 71.59 ;
      RECT 27.245 71.59 27.775 71.725 ;
      RECT 27.065 56.84 27.955 63.63 ;
      RECT 25.86 56.9 26.39 63.57 ;
      RECT 25.87 63.57 26.38 63.63 ;
      RECT 25.87 56.84 26.38 56.9 ;
      RECT 28.63 56.9 29.16 63.57 ;
      RECT 28.64 63.57 29.15 63.63 ;
      RECT 28.64 56.84 29.15 56.9 ;
      RECT 28.63 66.9 29.16 71.725 ;
      RECT 28.64 66.84 29.15 66.9 ;
      RECT 25.86 66.9 26.39 71.725 ;
      RECT 25.87 66.84 26.38 66.9 ;
      RECT 29.835 66.84 30.725 71.59 ;
      RECT 30.015 71.59 30.545 71.725 ;
      RECT 29.835 56.84 30.725 63.63 ;
      RECT 31.4 56.9 31.93 63.57 ;
      RECT 31.41 63.57 31.92 63.63 ;
      RECT 31.41 56.84 31.92 56.9 ;
      RECT 31.4 66.9 31.93 71.725 ;
      RECT 31.41 66.84 31.92 66.9 ;
      RECT 35.375 66.84 36.265 71.59 ;
      RECT 24.295 36.84 25.185 43.63 ;
      RECT 21.525 36.84 22.415 43.63 ;
      RECT 24.295 26.84 25.185 33.63 ;
      RECT 21.525 26.84 22.415 33.63 ;
      RECT 24.295 46.84 25.185 53.63 ;
      RECT 21.525 46.84 22.415 53.63 ;
      RECT 23.09 46.9 23.62 53.57 ;
      RECT 23.1 53.57 23.61 53.63 ;
      RECT 23.1 46.84 23.61 46.9 ;
      RECT 23.09 36.9 23.62 43.57 ;
      RECT 23.1 43.57 23.61 43.63 ;
      RECT 23.1 36.84 23.61 36.9 ;
      RECT 23.09 26.9 23.62 33.57 ;
      RECT 23.1 33.57 23.61 33.63 ;
      RECT 23.1 26.84 23.61 26.9 ;
      RECT 27.065 36.84 27.955 43.63 ;
      RECT 27.065 26.84 27.955 33.63 ;
      RECT 27.065 46.84 27.955 53.63 ;
      RECT 28.63 46.9 29.16 53.57 ;
      RECT 28.64 53.57 29.15 53.63 ;
      RECT 28.64 46.84 29.15 46.9 ;
      RECT 25.86 46.9 26.39 53.57 ;
      RECT 25.87 53.57 26.38 53.63 ;
      RECT 25.87 46.84 26.38 46.9 ;
      RECT 25.86 36.9 26.39 43.57 ;
      RECT 25.87 43.57 26.38 43.63 ;
      RECT 25.87 36.84 26.38 36.9 ;
      RECT 28.63 36.9 29.16 43.57 ;
      RECT 28.64 43.57 29.15 43.63 ;
      RECT 28.64 36.84 29.15 36.9 ;
      RECT 25.86 26.9 26.39 33.57 ;
      RECT 25.87 33.57 26.38 33.63 ;
      RECT 25.87 26.84 26.38 26.9 ;
      RECT 28.63 26.9 29.16 33.57 ;
      RECT 28.64 33.57 29.15 33.63 ;
      RECT 28.64 26.84 29.15 26.9 ;
      RECT 29.835 36.84 30.725 43.63 ;
      RECT 29.835 26.84 30.725 33.63 ;
      RECT 29.835 46.84 30.725 53.63 ;
      RECT 31.4 46.9 31.93 53.57 ;
      RECT 31.41 53.57 31.92 53.63 ;
      RECT 31.41 46.84 31.92 46.9 ;
      RECT 31.4 36.9 31.93 43.57 ;
      RECT 31.41 43.57 31.92 43.63 ;
      RECT 31.41 36.84 31.92 36.9 ;
      RECT 31.4 26.9 31.93 33.57 ;
      RECT 31.41 33.57 31.92 33.63 ;
      RECT 31.41 26.84 31.92 26.9 ;
      RECT 35.375 36.84 36.265 43.63 ;
      RECT 32.605 36.84 33.495 43.63 ;
      RECT 35.375 26.84 36.265 33.63 ;
      RECT 32.605 26.84 33.495 33.63 ;
      RECT 35.375 46.84 36.265 53.63 ;
      RECT 32.605 46.84 33.495 53.63 ;
      RECT 34.17 46.9 34.7 53.57 ;
      RECT 34.18 53.57 34.69 53.63 ;
      RECT 34.18 46.84 34.69 46.9 ;
      RECT 34.17 36.9 34.7 43.57 ;
      RECT 34.18 43.57 34.69 43.63 ;
      RECT 34.18 36.84 34.69 36.9 ;
      RECT 34.17 26.9 34.7 33.57 ;
      RECT 34.18 33.57 34.69 33.63 ;
      RECT 34.18 26.84 34.69 26.9 ;
      RECT 38.145 36.84 39.035 43.63 ;
      RECT 38.145 26.84 39.035 33.63 ;
      RECT 38.145 46.84 39.035 53.63 ;
      RECT 36.94 46.9 37.47 53.57 ;
      RECT 36.95 53.57 37.46 53.63 ;
      RECT 36.95 46.84 37.46 46.9 ;
      RECT 36.94 36.9 37.47 43.57 ;
      RECT 36.95 43.57 37.46 43.63 ;
      RECT 36.95 36.84 37.46 36.9 ;
      RECT 36.94 26.9 37.47 33.57 ;
      RECT 36.95 33.57 37.46 33.63 ;
      RECT 36.95 26.84 37.46 26.9 ;
      RECT 39.71 26.9 40.24 33.57 ;
      RECT 39.72 33.57 40.23 33.63 ;
      RECT 39.72 26.84 40.23 26.9 ;
      RECT 39.71 46.9 40.24 53.57 ;
      RECT 39.72 53.57 40.23 53.63 ;
      RECT 39.72 46.84 40.23 46.9 ;
      RECT 39.71 36.9 40.24 43.57 ;
      RECT 39.72 43.57 40.23 43.63 ;
      RECT 39.72 36.84 40.23 36.9 ;
      RECT 43.685 36.84 44.575 43.63 ;
      RECT 40.915 36.84 41.805 43.63 ;
      RECT 43.685 26.84 44.575 33.63 ;
      RECT 40.915 26.84 41.805 33.63 ;
      RECT 43.685 46.84 44.575 53.63 ;
      RECT 40.915 46.84 41.805 53.63 ;
      RECT 42.48 26.9 43.01 33.57 ;
      RECT 42.49 33.57 43 33.63 ;
      RECT 42.49 26.84 43 26.9 ;
      RECT 42.48 46.9 43.01 53.57 ;
      RECT 42.49 53.57 43 53.63 ;
      RECT 42.49 46.84 43 46.9 ;
      RECT 42.48 36.9 43.01 43.57 ;
      RECT 42.49 43.57 43 43.63 ;
      RECT 42.49 36.84 43 36.9 ;
      RECT 46.455 36.84 47.345 43.63 ;
      RECT 46.455 26.84 47.345 33.63 ;
      RECT 46.455 46.84 47.345 53.63 ;
      RECT 45.25 26.9 45.78 33.57 ;
      RECT 45.26 33.57 45.77 33.63 ;
      RECT 45.26 26.84 45.77 26.9 ;
      RECT 45.25 46.9 45.78 53.57 ;
      RECT 45.26 53.57 45.77 53.63 ;
      RECT 45.26 46.84 45.77 46.9 ;
      RECT 45.25 36.9 45.78 43.57 ;
      RECT 45.26 43.57 45.77 43.63 ;
      RECT 45.26 36.84 45.77 36.9 ;
      RECT 49.225 36.84 50.115 43.63 ;
      RECT 49.225 26.84 50.115 33.63 ;
      RECT 49.225 46.84 50.115 53.63 ;
      RECT 48.02 26.9 48.55 33.57 ;
      RECT 48.03 33.57 48.54 33.63 ;
      RECT 48.03 26.84 48.54 26.9 ;
      RECT 50.79 26.9 51.32 33.57 ;
      RECT 50.8 33.57 51.31 33.63 ;
      RECT 50.8 26.84 51.31 26.9 ;
      RECT 48.02 46.9 48.55 53.57 ;
      RECT 48.03 53.57 48.54 53.63 ;
      RECT 48.03 46.84 48.54 46.9 ;
      RECT 50.79 46.9 51.32 53.57 ;
      RECT 50.8 53.57 51.31 53.63 ;
      RECT 50.8 46.84 51.31 46.9 ;
      RECT 48.02 36.9 48.55 43.57 ;
      RECT 1.84 17.21 2.995 18.69 ;
      RECT 1.35 17.04 7.11 17.21 ;
      RECT 6.94 1.19 7.11 17.04 ;
      RECT 1.35 1.02 7.11 1.19 ;
      RECT 0.24 18.69 2.995 19.2 ;
      RECT 1.35 1.19 1.52 17.04 ;
      RECT 1.845 9.65 2.015 16.61 ;
      RECT 1.845 2 2.015 8.96 ;
      RECT 1.76 20.14 2.685 23.06 ;
      RECT 1.76 19.63 9.385 20.14 ;
      RECT 5.525 9.65 5.695 16.61 ;
      RECT 5.525 2 5.695 8.96 ;
      RECT 5.065 9.65 5.235 16.44 ;
      RECT 5.065 2 5.235 8.96 ;
      RECT 4.605 9.65 4.775 16.61 ;
      RECT 4.605 2 4.775 8.96 ;
      RECT 4.145 9.65 4.315 16.44 ;
      RECT 4.145 2 4.315 8.96 ;
      RECT 3.685 9.65 3.855 16.61 ;
      RECT 3.685 2 3.855 8.96 ;
      RECT 3.225 9.65 3.395 16.44 ;
      RECT 3.225 2 3.395 8.96 ;
      RECT 2.765 9.65 2.935 16.61 ;
      RECT 2.765 2 2.935 8.96 ;
      RECT 2.305 9.65 2.475 16.44 ;
      RECT 2.305 2 2.475 8.96 ;
      RECT 5.89 23.01 10.65 23.015 ;
      RECT 4.975 22.29 10.65 23.01 ;
      RECT 5.985 9.65 6.155 16.44 ;
      RECT 5.985 2 6.155 8.96 ;
      RECT 6.445 9.65 6.615 16.61 ;
      RECT 6.445 2 6.615 8.96 ;
      RECT 56.155 1.28 56.565 17.04 ;
      RECT 8.345 17.58 16.645 18.35 ;
      RECT 36.165 1.28 37.055 17.04 ;
      RECT 16.655 0.51 56.565 1.28 ;
      RECT 16.655 1.28 17.065 1.41 ;
      RECT 8.345 17.45 16.655 17.58 ;
      RECT 8.345 17.04 56.565 17.45 ;
      RECT 8.345 1.41 17.065 17.04 ;
      RECT 17.625 1.48 19.125 16.48 ;
      RECT 19.685 1.48 21.185 16.48 ;
      RECT 21.745 1.48 23.245 16.48 ;
      RECT 23.805 1.48 25.305 16.48 ;
      RECT 25.865 1.48 27.365 16.48 ;
      RECT 27.925 1.48 29.425 16.48 ;
      RECT 29.985 1.48 31.485 16.48 ;
      RECT 32.045 1.48 33.545 16.48 ;
      RECT 34.105 1.48 35.605 16.48 ;
      RECT 37.615 1.48 39.115 16.48 ;
      RECT 39.675 1.48 41.175 16.48 ;
      RECT 41.735 1.48 43.235 16.48 ;
      RECT 43.795 1.48 45.295 16.48 ;
      RECT 45.855 1.48 47.355 16.48 ;
      RECT 47.915 1.48 49.415 16.48 ;
      RECT 49.975 1.48 51.475 16.48 ;
      RECT 54.095 1.48 55.595 16.48 ;
      RECT 52.035 1.48 53.535 16.48 ;
      RECT 56.98 16.365 57.51 16.895 ;
      RECT 66.7 1.205 67.23 1.735 ;
      RECT 66.785 1.735 67.115 1.745 ;
      RECT 69.53 19.01 70.265 19.61 ;
      RECT 70.495 17.96 71.095 18.695 ;
      RECT 70.87 2.06 71.04 9.02 ;
      RECT 70.87 9.71 71.04 16.67 ;
      RECT 70.41 2.06 70.58 9.02 ;
      RECT 70.41 9.71 70.58 16.5 ;
      RECT 69.95 2.06 70.12 9.02 ;
      RECT 69.95 9.71 70.12 16.67 ;
      RECT 69.49 2.06 69.66 9.02 ;
      RECT 69.49 9.71 69.66 16.5 ;
      RECT 69.03 2.06 69.2 9.02 ;
      RECT 69.03 9.71 69.2 16.67 ;
      RECT 68.57 2.06 68.74 9.02 ;
      RECT 68.57 9.71 68.74 16.5 ;
      RECT 68.11 2.06 68.28 9.02 ;
      RECT 68.11 9.71 68.28 16.67 ;
      RECT 67.615 17.1 73.375 17.27 ;
      RECT 73.205 1.25 73.375 17.1 ;
      RECT 67.61 1.08 73.375 1.25 ;
      RECT 67.615 1.25 67.785 17.1 ;
      RECT 72.25 9.71 72.42 16.5 ;
      RECT 71.79 2.06 71.96 9.02 ;
      RECT 71.79 9.71 71.96 16.67 ;
      RECT 71.33 2.06 71.5 9.02 ;
      RECT 71.33 9.71 71.5 16.5 ;
      RECT 72.71 2.06 72.88 9.02 ;
      RECT 72.71 9.71 72.88 16.67 ;
      RECT 72.25 2.06 72.42 9.02 ;
      RECT 13.215 36.84 14.105 43.63 ;
      RECT 13.215 26.84 14.105 33.63 ;
      RECT 13.215 46.84 14.105 53.63 ;
      RECT 13.06 44.1 65.59 46.62 ;
      RECT 13.19 34.1 65.59 36.62 ;
      RECT 15.985 36.84 16.875 43.63 ;
      RECT 15.985 26.84 16.875 33.63 ;
      RECT 15.985 46.84 16.875 53.63 ;
      RECT 14.78 26.9 15.31 33.57 ;
      RECT 14.79 33.57 15.3 33.63 ;
      RECT 14.79 26.84 15.3 26.9 ;
      RECT 14.78 36.9 15.31 43.57 ;
      RECT 14.79 43.57 15.3 43.63 ;
      RECT 14.79 36.84 15.3 36.9 ;
      RECT 14.78 46.9 15.31 53.57 ;
      RECT 14.79 53.57 15.3 53.63 ;
      RECT 14.79 46.84 15.3 46.9 ;
      RECT 18.755 36.84 19.645 43.63 ;
      RECT 18.755 26.84 19.645 33.63 ;
      RECT 18.755 46.84 19.645 53.63 ;
      RECT 17.55 36.9 18.08 43.57 ;
      RECT 17.56 43.57 18.07 43.63 ;
      RECT 17.56 36.84 18.07 36.9 ;
      RECT 20.32 36.9 20.85 43.57 ;
      RECT 20.33 43.57 20.84 43.63 ;
      RECT 20.33 36.84 20.84 36.9 ;
      RECT 17.55 26.9 18.08 33.57 ;
      RECT 17.56 33.57 18.07 33.63 ;
      RECT 17.56 26.84 18.07 26.9 ;
      RECT 20.32 26.9 20.85 33.57 ;
      RECT 20.33 33.57 20.84 33.63 ;
      RECT 20.33 26.84 20.84 26.9 ;
      RECT 17.55 46.9 18.08 53.57 ;
      RECT 17.56 53.57 18.07 53.63 ;
      RECT 17.56 46.84 18.07 46.9 ;
      RECT 20.32 46.9 20.85 53.57 ;
      RECT 20.33 53.57 20.84 53.63 ;
      RECT 20.33 46.84 20.84 46.9 ;
      RECT 21.57 83.15 21.74 99.925 ;
      RECT 9.69 23.825 69.72 24.355 ;
      RECT 9.155 197.35 69.72 197.38 ;
      RECT 8.975 196.85 69.72 197.35 ;
      RECT 9.675 98.165 10.28 99.49 ;
      RECT 9.69 82.98 21.74 83.15 ;
      RECT 69.19 100.095 69.72 196.85 ;
      RECT 21.57 99.925 69.72 100.095 ;
      RECT 69.19 24.355 69.72 99.925 ;
      RECT 9.73 99.49 10.28 106.965 ;
      RECT 8.975 144.535 10.28 196.85 ;
      RECT 9.155 106.965 10.28 144.535 ;
      RECT 9.69 83.15 10.28 98.165 ;
      RECT 9.69 24.355 10.28 82.98 ;
      RECT 22.77 98.99 68.14 99.16 ;
      RECT 12 82.21 12.505 82.255 ;
      RECT 12.455 81.7 23.28 81.745 ;
      RECT 11.37 43.62 12.22 46.905 ;
      RECT 67.29 26.085 68.14 82.18 ;
      RECT 22.43 90.845 23.28 97.89 ;
      RECT 22.43 82.35 23.28 90.675 ;
      RECT 22.77 97.89 23.28 98.99 ;
      RECT 67.29 90.845 68.14 98.99 ;
      RECT 22.43 90.675 68.14 90.845 ;
      RECT 67.29 82.35 68.14 90.675 ;
      RECT 11.275 26.085 12.22 34.04 ;
      RECT 11.37 34.04 12.22 36.745 ;
      RECT 11.37 81.435 12.22 81.745 ;
      RECT 11.37 81.745 23.28 82.18 ;
      RECT 22.43 82.21 68.14 82.35 ;
      RECT 11.37 82.18 68.14 82.21 ;
      RECT 11.275 36.745 12.22 43.62 ;
      RECT 11.275 25.065 68.14 26.085 ;
      RECT 11.275 46.905 12.22 81.435 ;
      RECT 11.04 144.465 21.49 145.315 ;
      RECT 11.04 194.935 68.495 195.885 ;
      RECT 20.64 100.865 68.495 101.035 ;
      RECT 20.64 117.94 21.49 144.465 ;
      RECT 67.575 100.84 68.495 100.865 ;
      RECT 20.64 109.445 21.49 117.77 ;
      RECT 20.64 101.035 21.49 109.275 ;
      RECT 20.64 109.275 68.495 109.445 ;
      RECT 67.575 117.94 68.495 194.935 ;
      RECT 20.64 117.77 68.495 117.94 ;
      RECT 67.575 109.445 68.495 117.77 ;
      RECT 67.575 101.035 68.495 109.275 ;
      RECT 11.04 145.315 12.22 194.935 ;
    LAYER met3 ;
      RECT 49.655 0 75 69.89 ;
      RECT 46.96 74.34 75 76.65 ;
      RECT 37.28 69.89 75 70.94 ;
      RECT 37.28 70.94 75 74.34 ;
      RECT 49.27 76.65 75 84.645 ;
      RECT 49.27 84.645 75 86.795 ;
      RECT 51.42 86.795 75 88.21 ;
      RECT 0 189.915 75 198 ;
      RECT 51.42 88.21 75 97.52 ;
      RECT 49.235 100.33 53.93 164.295 ;
      RECT 49.235 164.295 49.47 168.755 ;
      RECT 49.235 96.645 53.93 100.33 ;
      RECT 60.73 97.52 75 189.915 ;
      RECT 0 94.145 15.205 189.915 ;
      RECT 0 85.9 15.205 94.145 ;
      RECT 0 84.485 23.45 85.9 ;
      RECT 0 0 24.74 24.685 ;
      RECT 0 82.335 23.45 84.485 ;
      RECT 0 24.685 25.6 82.335 ;
      RECT 25.515 170.445 25.635 189.915 ;
      RECT 22.005 166.935 25.635 170.445 ;
      RECT 22.005 96.955 25.635 166.935 ;
      RECT 24.625 94.335 25.635 96.955 ;
      RECT 32.545 84.855 34.105 85.865 ;
      RECT 32.545 85.865 33.555 86.415 ;
      RECT 33.02 84.38 34.105 84.855 ;
      RECT 37.325 168.86 37.545 189.915 ;
      RECT 37.28 0 37.98 69.89 ;
      RECT 37.325 167.295 37.545 168.86 ;
      RECT 35.215 90.775 40.41 93.555 ;
      RECT 39.785 87.195 41.21 87.61 ;
      RECT 40.26 84.38 41.21 84.855 ;
      RECT 39.785 84.855 41.21 87.195 ;
      RECT 32.435 162.405 42.435 163.97 ;
      RECT 34 163.97 39.11 167.295 ;
      RECT 32.435 93.555 42.435 95.58 ;
      RECT 32.435 95.58 42.435 162.405 ;
      RECT 40.2 87.61 50.245 96.645 ;
      RECT 49.235 168.755 49.47 189.915 ;
      RECT 3.0 88.255 16.7 88.405 ;
      RECT 3.0 88.405 16.545 88.555 ;
      RECT 3.0 88.555 16.4 88.705 ;
      RECT 3.0 88.705 16.25 88.855 ;
      RECT 3.0 88.855 16.095 89.005 ;
      RECT 3.0 89.005 15.95 89.155 ;
      RECT 3.0 89.155 15.8 89.305 ;
      RECT 3.0 89.305 15.65 89.455 ;
      RECT 3.0 89.455 15.5 89.605 ;
      RECT 3.0 89.605 15.35 89.755 ;
      RECT 3.0 89.755 15.2 89.905 ;
      RECT 3.0 89.905 15.05 90.055 ;
      RECT 3.0 90.055 14.9 90.205 ;
      RECT 3.0 90.205 14.75 90.355 ;
      RECT 3.0 90.355 14.6 90.505 ;
      RECT 3.0 90.505 14.45 90.655 ;
      RECT 3.0 90.655 14.3 90.805 ;
      RECT 3.0 90.805 14.15 90.955 ;
      RECT 3.0 90.955 14.0 91.105 ;
      RECT 3.0 91.105 13.85 91.255 ;
      RECT 3.0 91.255 13.7 91.405 ;
      RECT 3.0 91.405 13.55 91.555 ;
      RECT 3.0 91.555 13.4 91.705 ;
      RECT 3.0 91.705 13.25 91.855 ;
      RECT 3.0 91.855 13.1 92.005 ;
      RECT 3.0 92.005 12.95 92.155 ;
      RECT 3.0 92.155 12.8 92.305 ;
      RECT 3.0 92.305 12.65 92.455 ;
      RECT 3.0 92.455 12.5 92.605 ;
      RECT 3.0 92.605 12.35 92.755 ;
      RECT 3.0 92.755 12.205 92.9 ;
      RECT 52.42 83.4 72.0 83.55 ;
      RECT 52.57 83.55 72.0 83.7 ;
      RECT 52.72 83.7 72.0 83.85 ;
      RECT 52.87 83.85 72.0 84 ;
      RECT 53.02 84 72.0 84.15 ;
      RECT 53.17 84.15 72.0 84.3 ;
      RECT 53.32 84.3 72.0 84.45 ;
      RECT 53.47 84.45 72.0 84.6 ;
      RECT 53.62 84.6 72.0 84.75 ;
      RECT 53.77 84.75 72.0 84.9 ;
      RECT 53.92 84.9 72.0 85.05 ;
      RECT 54.07 85.05 72.0 85.2 ;
      RECT 54.22 85.2 72.0 85.35 ;
      RECT 54.37 85.35 72.0 85.5 ;
      RECT 54.42 85.5 72.0 85.55 ;
      RECT 54.57 86.965 72.0 87.115 ;
      RECT 54.72 87.115 72.0 87.265 ;
      RECT 54.87 87.265 72.0 87.415 ;
      RECT 55.02 87.415 72.0 87.565 ;
      RECT 55.17 87.565 72.0 87.715 ;
      RECT 55.32 87.715 72.0 87.865 ;
      RECT 55.47 87.865 72.0 88.015 ;
      RECT 55.62 88.015 72.0 88.165 ;
      RECT 55.77 88.165 72.0 88.315 ;
      RECT 55.92 88.315 72.0 88.465 ;
      RECT 56.07 88.465 72.0 88.615 ;
      RECT 56.22 88.615 72.0 88.765 ;
      RECT 56.37 88.765 72.0 88.915 ;
      RECT 56.52 88.915 72.0 89.065 ;
      RECT 56.67 89.065 72.0 89.215 ;
      RECT 56.82 89.215 72.0 89.365 ;
      RECT 56.97 89.365 72.0 89.515 ;
      RECT 57.12 89.515 72.0 89.665 ;
      RECT 57.27 89.665 72.0 89.815 ;
      RECT 57.42 89.815 72.0 89.965 ;
      RECT 57.57 89.965 72.0 90.115 ;
      RECT 57.72 90.115 72.0 90.265 ;
      RECT 57.87 90.265 72.0 90.415 ;
      RECT 58.02 90.415 72.0 90.565 ;
      RECT 58.17 90.565 72.0 90.715 ;
      RECT 58.32 90.715 72.0 90.865 ;
      RECT 58.47 90.865 72.0 91.015 ;
      RECT 58.62 91.015 72.0 91.165 ;
      RECT 58.77 91.165 72.0 91.315 ;
      RECT 58.92 91.315 72.0 91.465 ;
      RECT 59.07 91.465 72.0 91.615 ;
      RECT 59.22 91.615 72.0 91.765 ;
      RECT 59.37 91.765 72.0 91.915 ;
      RECT 59.52 91.915 72.0 92.065 ;
      RECT 59.67 92.065 72.0 92.215 ;
      RECT 59.82 92.215 72.0 92.365 ;
      RECT 59.97 92.365 72.0 92.515 ;
      RECT 60.12 92.515 72.0 92.665 ;
      RECT 60.27 92.665 72.0 92.815 ;
      RECT 60.42 92.815 72.0 92.965 ;
      RECT 60.57 92.965 72.0 93.115 ;
      RECT 60.72 93.115 72.0 93.265 ;
      RECT 60.87 93.265 72.0 93.415 ;
      RECT 61.02 93.415 72.0 93.565 ;
      RECT 61.17 93.565 72.0 93.715 ;
      RECT 61.32 93.715 72.0 93.865 ;
      RECT 61.47 93.865 72.0 94.015 ;
      RECT 61.62 94.015 72.0 94.165 ;
      RECT 61.77 94.165 72.0 94.315 ;
      RECT 61.92 94.315 72.0 94.465 ;
      RECT 62.07 94.465 72.0 94.615 ;
      RECT 62.22 94.615 72.0 94.765 ;
      RECT 62.37 94.765 72.0 94.915 ;
      RECT 62.52 94.915 72.0 95.065 ;
      RECT 62.67 95.065 72.0 95.215 ;
      RECT 62.82 95.215 72.0 95.365 ;
      RECT 62.97 95.365 72.0 95.515 ;
      RECT 63.12 95.515 72.0 95.665 ;
      RECT 63.27 95.665 72.0 95.815 ;
      RECT 63.42 95.815 72.0 95.965 ;
      RECT 63.57 95.965 72.0 96.115 ;
      RECT 63.72 96.115 72.0 96.265 ;
      RECT 63.73 96.265 72.0 96.275 ;
      RECT 49.905 72.89 72.0 73.04 ;
      RECT 50.055 73.04 72.0 73.19 ;
      RECT 50.205 73.19 72.0 73.34 ;
      RECT 50.355 73.34 72.0 73.49 ;
      RECT 50.505 73.49 72.0 73.64 ;
      RECT 50.655 73.64 72.0 73.79 ;
      RECT 50.805 73.79 72.0 73.94 ;
      RECT 50.955 73.94 72.0 74.09 ;
      RECT 51.105 74.09 72.0 74.24 ;
      RECT 51.255 74.24 72.0 74.39 ;
      RECT 51.405 74.39 72.0 74.54 ;
      RECT 51.555 74.54 72.0 74.69 ;
      RECT 51.705 74.69 72.0 74.84 ;
      RECT 51.855 74.84 72.0 74.99 ;
      RECT 52.005 74.99 72.0 75.14 ;
      RECT 52.155 75.14 72.0 75.29 ;
      RECT 52.27 75.29 72.0 75.405 ;
      RECT 53.62 84.6 72.0 84.75 ;
      RECT 53.77 84.75 72.0 84.9 ;
      RECT 53.92 84.9 72.0 85.05 ;
      RECT 54.07 85.05 72.0 85.2 ;
      RECT 54.22 85.2 72.0 85.35 ;
      RECT 54.37 85.35 72.0 85.5 ;
      RECT 54.42 85.5 72.0 85.55 ;
      RECT 54.57 86.965 72.0 87.115 ;
      RECT 54.72 87.115 72.0 87.265 ;
      RECT 54.87 87.265 72.0 87.415 ;
      RECT 55.02 87.415 72.0 87.565 ;
      RECT 55.17 87.565 72.0 87.715 ;
      RECT 55.32 87.715 72.0 87.865 ;
      RECT 55.47 87.865 72.0 88.015 ;
      RECT 55.62 88.015 72.0 88.165 ;
      RECT 55.77 88.165 72.0 88.315 ;
      RECT 55.92 88.315 72.0 88.465 ;
      RECT 56.07 88.465 72.0 88.615 ;
      RECT 56.22 88.615 72.0 88.765 ;
      RECT 56.37 88.765 72.0 88.915 ;
      RECT 56.52 88.915 72.0 89.065 ;
      RECT 56.67 89.065 72.0 89.215 ;
      RECT 56.82 89.215 72.0 89.365 ;
      RECT 56.97 89.365 72.0 89.515 ;
      RECT 57.12 89.515 72.0 89.665 ;
      RECT 57.27 89.665 72.0 89.815 ;
      RECT 57.42 89.815 72.0 89.965 ;
      RECT 57.57 89.965 72.0 90.115 ;
      RECT 57.72 90.115 72.0 90.265 ;
      RECT 57.87 90.265 72.0 90.415 ;
      RECT 58.02 90.415 72.0 90.565 ;
      RECT 58.17 90.565 72.0 90.715 ;
      RECT 58.32 90.715 72.0 90.865 ;
      RECT 58.47 90.865 72.0 91.015 ;
      RECT 58.62 91.015 72.0 91.165 ;
      RECT 58.77 91.165 72.0 91.315 ;
      RECT 58.92 91.315 72.0 91.465 ;
      RECT 59.07 91.465 72.0 91.615 ;
      RECT 59.22 91.615 72.0 91.765 ;
      RECT 59.37 91.765 72.0 91.915 ;
      RECT 59.52 91.915 72.0 92.065 ;
      RECT 59.67 92.065 72.0 92.215 ;
      RECT 59.82 92.215 72.0 92.365 ;
      RECT 59.97 92.365 72.0 92.515 ;
      RECT 60.12 92.515 72.0 92.665 ;
      RECT 60.27 92.665 72.0 92.815 ;
      RECT 60.42 92.815 72.0 92.965 ;
      RECT 60.57 92.965 72.0 93.115 ;
      RECT 60.72 93.115 72.0 93.265 ;
      RECT 60.87 93.265 72.0 93.415 ;
      RECT 61.02 93.415 72.0 93.565 ;
      RECT 61.17 93.565 72.0 93.715 ;
      RECT 61.32 93.715 72.0 93.865 ;
      RECT 61.47 93.865 72.0 94.015 ;
      RECT 61.62 94.015 72.0 94.165 ;
      RECT 61.77 94.165 72.0 94.315 ;
      RECT 61.92 94.315 72.0 94.465 ;
      RECT 62.07 94.465 72.0 94.615 ;
      RECT 62.22 94.615 72.0 94.765 ;
      RECT 62.37 94.765 72.0 94.915 ;
      RECT 62.52 94.915 72.0 95.065 ;
      RECT 62.67 95.065 72.0 95.215 ;
      RECT 62.82 95.215 72.0 95.365 ;
      RECT 62.97 95.365 72.0 95.515 ;
      RECT 63.12 95.515 72.0 95.665 ;
      RECT 63.27 95.665 72.0 95.815 ;
      RECT 63.42 95.815 72.0 95.965 ;
      RECT 63.57 95.965 72.0 96.115 ;
      RECT 63.72 96.115 72.0 96.265 ;
      RECT 63.73 96.265 72.0 96.275 ;
      RECT 20.45 84.655 23.45 84.805 ;
      RECT 20.295 84.805 23.45 84.955 ;
      RECT 20.15 84.955 23.45 85.105 ;
      RECT 20.0 85.105 23.45 85.255 ;
      RECT 19.845 85.255 23.45 85.405 ;
      RECT 19.7 85.405 23.45 85.555 ;
      RECT 19.545 85.555 23.45 85.705 ;
      RECT 19.4 85.705 23.45 85.855 ;
      RECT 19.25 85.855 23.45 85.9 ;
      RECT 51.42 86.965 54.42 87.115 ;
      RECT 51.42 87.115 54.57 87.265 ;
      RECT 51.42 87.265 54.72 87.415 ;
      RECT 51.42 87.415 54.87 87.565 ;
      RECT 51.42 87.565 55.02 87.715 ;
      RECT 51.42 87.715 55.17 87.865 ;
      RECT 51.42 87.865 55.32 88.015 ;
      RECT 51.42 88.015 55.47 88.165 ;
      RECT 51.42 88.165 55.62 88.21 ;
      RECT 3.0 81.09 22.45 81.24 ;
      RECT 3.0 81.24 22.295 81.39 ;
      RECT 3.0 81.39 22.15 81.54 ;
      RECT 3.0 81.54 22.0 81.69 ;
      RECT 3.0 81.69 21.845 81.84 ;
      RECT 3.0 81.84 21.7 81.99 ;
      RECT 3.0 81.99 21.545 82.14 ;
      RECT 3.0 82.14 21.4 82.29 ;
      RECT 3.0 82.29 21.25 82.44 ;
      RECT 3.0 82.44 21.095 82.59 ;
      RECT 3.0 82.59 20.95 82.74 ;
      RECT 3.0 82.74 20.795 82.89 ;
      RECT 3.0 82.89 20.65 83.04 ;
      RECT 3.0 83.04 20.5 83.19 ;
      RECT 3.0 83.19 20.45 83.24 ;
      RECT 3.0 84.655 20.295 84.805 ;
      RECT 3.0 84.805 20.15 84.955 ;
      RECT 3.0 84.955 20.0 85.105 ;
      RECT 3.0 85.105 19.845 85.255 ;
      RECT 3.0 85.255 19.7 85.405 ;
      RECT 3.0 85.405 19.545 85.555 ;
      RECT 3.0 85.555 19.4 85.705 ;
      RECT 3.0 85.705 19.25 85.855 ;
      RECT 3.0 85.855 19.095 86.005 ;
      RECT 3.0 86.005 18.95 86.155 ;
      RECT 3.0 86.155 18.795 86.305 ;
      RECT 3.0 86.305 18.65 86.455 ;
      RECT 3.0 86.455 18.5 86.605 ;
      RECT 3.0 86.605 18.345 86.755 ;
      RECT 3.0 86.755 18.2 86.905 ;
      RECT 3.0 86.905 18.045 87.055 ;
      RECT 3.0 87.055 17.9 87.205 ;
      RECT 3.0 87.205 17.75 87.355 ;
      RECT 3.0 87.355 17.595 87.505 ;
      RECT 3.0 87.505 17.45 87.655 ;
      RECT 3.0 87.655 17.295 87.805 ;
      RECT 3.0 87.805 17.15 87.955 ;
      RECT 3.0 87.955 17.0 88.105 ;
      RECT 3.0 88.105 16.845 88.255 ;
      RECT 56.22 92.86 75 93.01 ;
      RECT 56.37 93.01 75 93.16 ;
      RECT 56.52 93.16 75 93.31 ;
      RECT 56.67 93.31 75 93.46 ;
      RECT 56.82 93.46 75 93.61 ;
      RECT 56.97 93.61 75 93.76 ;
      RECT 57.12 93.76 75 93.91 ;
      RECT 57.27 93.91 75 94.06 ;
      RECT 57.42 94.06 75 94.21 ;
      RECT 57.57 94.21 75 94.36 ;
      RECT 57.72 94.36 75 94.51 ;
      RECT 57.87 94.51 75 94.66 ;
      RECT 58.02 94.66 75 94.81 ;
      RECT 58.17 94.81 75 94.96 ;
      RECT 58.32 94.96 75 95.11 ;
      RECT 58.47 95.11 75 95.26 ;
      RECT 58.62 95.26 75 95.41 ;
      RECT 58.77 95.41 75 95.56 ;
      RECT 58.92 95.56 75 95.71 ;
      RECT 59.07 95.71 75 95.86 ;
      RECT 59.22 95.86 75 96.01 ;
      RECT 59.37 96.01 75 96.16 ;
      RECT 59.52 96.16 75 96.31 ;
      RECT 59.67 96.31 75 96.46 ;
      RECT 59.82 96.46 75 96.61 ;
      RECT 59.97 96.61 75 96.76 ;
      RECT 60.12 96.76 75 96.91 ;
      RECT 60.27 96.91 75 97.06 ;
      RECT 60.42 97.06 75 97.21 ;
      RECT 60.57 97.21 75 97.36 ;
      RECT 60.72 97.36 75 97.51 ;
      RECT 60.73 97.51 75 97.52 ;
      RECT 3.0 81.09 22.45 81.24 ;
      RECT 3.0 81.24 22.295 81.39 ;
      RECT 3.0 81.39 22.15 81.54 ;
      RECT 3.0 81.54 22.0 81.69 ;
      RECT 3.0 81.69 21.845 81.84 ;
      RECT 3.0 81.84 21.7 81.99 ;
      RECT 3.0 81.99 21.545 82.14 ;
      RECT 3.0 82.14 21.4 82.29 ;
      RECT 3.0 82.29 21.25 82.44 ;
      RECT 3.0 82.44 21.095 82.59 ;
      RECT 3.0 82.59 20.95 82.74 ;
      RECT 3.0 82.74 20.795 82.89 ;
      RECT 3.0 82.89 20.65 83.04 ;
      RECT 3.0 83.04 20.5 83.19 ;
      RECT 3.0 83.19 20.45 83.24 ;
      RECT 3.0 84.655 20.295 84.805 ;
      RECT 3.0 84.805 20.15 84.955 ;
      RECT 3.0 84.955 20.0 85.105 ;
      RECT 3.0 85.105 19.845 85.255 ;
      RECT 3.0 85.255 19.7 85.405 ;
      RECT 3.0 85.405 19.545 85.555 ;
      RECT 3.0 85.555 19.4 85.705 ;
      RECT 3.0 85.705 19.25 85.855 ;
      RECT 3.0 85.855 19.095 86.005 ;
      RECT 3.0 86.005 18.95 86.155 ;
      RECT 3.0 86.155 18.795 86.305 ;
      RECT 3.0 86.305 18.65 86.455 ;
      RECT 3.0 86.455 18.5 86.605 ;
      RECT 3.0 86.605 18.345 86.755 ;
      RECT 3.0 86.755 18.2 86.905 ;
      RECT 3.0 86.905 18.045 87.055 ;
      RECT 3.0 87.055 17.9 87.205 ;
      RECT 3.0 87.205 17.75 87.355 ;
      RECT 3.0 87.355 17.595 87.505 ;
      RECT 3.0 87.505 17.45 87.655 ;
      RECT 3.0 87.655 17.295 87.805 ;
      RECT 3.0 87.805 17.15 87.955 ;
      RECT 3.0 87.955 17.0 88.105 ;
      RECT 3.0 88.105 16.845 88.255 ;
      RECT 3.0 88.255 16.7 88.405 ;
      RECT 3.0 88.405 16.545 88.555 ;
      RECT 3.0 88.555 16.4 88.705 ;
      RECT 3.0 88.705 16.25 88.855 ;
      RECT 3.0 88.855 16.095 89.005 ;
      RECT 3.0 89.005 15.95 89.155 ;
      RECT 3.0 89.155 15.8 89.305 ;
      RECT 3.0 89.305 15.65 89.455 ;
      RECT 3.0 89.455 15.5 89.605 ;
      RECT 3.0 89.605 15.35 89.755 ;
      RECT 3.0 89.755 15.2 89.905 ;
      RECT 3.0 89.905 15.05 90.055 ;
      RECT 3.0 90.055 14.9 90.205 ;
      RECT 3.0 90.205 14.75 90.355 ;
      RECT 3.0 90.355 14.6 90.505 ;
      RECT 3.0 90.505 14.45 90.655 ;
      RECT 3.0 90.655 14.3 90.805 ;
      RECT 3.0 90.805 14.15 90.955 ;
      RECT 3.0 90.955 14.0 91.105 ;
      RECT 3.0 91.105 13.85 91.255 ;
      RECT 3.0 91.255 13.7 91.405 ;
      RECT 3.0 91.405 13.55 91.555 ;
      RECT 3.0 91.555 13.4 91.705 ;
      RECT 3.0 91.705 13.25 91.855 ;
      RECT 3.0 91.855 13.1 92.005 ;
      RECT 3.0 92.005 12.95 92.155 ;
      RECT 3.0 92.155 12.8 92.305 ;
      RECT 3.0 92.305 12.65 92.455 ;
      RECT 3.0 92.455 12.5 92.605 ;
      RECT 3.0 92.605 12.35 92.755 ;
      RECT 3.0 92.755 12.205 92.9 ;
      RECT 49.905 72.89 72.0 73.04 ;
      RECT 50.055 73.04 72.0 73.19 ;
      RECT 50.205 73.19 72.0 73.34 ;
      RECT 50.355 73.34 72.0 73.49 ;
      RECT 50.505 73.49 72.0 73.64 ;
      RECT 50.655 73.64 72.0 73.79 ;
      RECT 50.805 73.79 72.0 73.94 ;
      RECT 50.955 73.94 72.0 74.09 ;
      RECT 51.105 74.09 72.0 74.24 ;
      RECT 51.255 74.24 72.0 74.39 ;
      RECT 51.405 74.39 72.0 74.54 ;
      RECT 51.555 74.54 72.0 74.69 ;
      RECT 51.705 74.69 72.0 74.84 ;
      RECT 51.855 74.84 72.0 74.99 ;
      RECT 52.005 74.99 72.0 75.14 ;
      RECT 52.155 75.14 72.0 75.29 ;
      RECT 52.27 75.29 72.0 75.405 ;
      RECT 52.42 83.4 72.0 83.55 ;
      RECT 52.57 83.55 72.0 83.7 ;
      RECT 52.72 83.7 72.0 83.85 ;
      RECT 52.87 83.85 72.0 84 ;
      RECT 53.02 84 72.0 84.15 ;
      RECT 53.17 84.15 72.0 84.3 ;
      RECT 53.32 84.3 72.0 84.45 ;
      RECT 53.47 84.45 72.0 84.6 ;
      RECT 48.45 95.71 49.31 95.86 ;
      RECT 48.6 95.86 49.46 96.01 ;
      RECT 48.75 96.01 49.61 96.16 ;
      RECT 48.9 96.16 49.76 96.31 ;
      RECT 49.05 96.31 49.91 96.46 ;
      RECT 49.2 96.46 50.06 96.61 ;
      RECT 49.235 96.61 50.21 96.645 ;
      RECT 47.11 74.34 75 74.49 ;
      RECT 47.26 74.49 75 74.64 ;
      RECT 47.41 74.64 75 74.79 ;
      RECT 47.56 74.79 75 74.94 ;
      RECT 47.71 74.94 75 75.09 ;
      RECT 47.86 75.09 75 75.24 ;
      RECT 48.01 75.24 75 75.39 ;
      RECT 48.16 75.39 75 75.54 ;
      RECT 48.31 75.54 75 75.69 ;
      RECT 48.46 75.69 75 75.84 ;
      RECT 48.61 75.84 75 75.99 ;
      RECT 48.76 75.99 75 76.14 ;
      RECT 48.91 76.14 75 76.29 ;
      RECT 49.06 76.29 75 76.44 ;
      RECT 49.21 76.44 75 76.59 ;
      RECT 49.27 76.59 75 76.65 ;
      RECT 49.235 96.645 50.245 96.795 ;
      RECT 49.235 96.795 50.395 96.945 ;
      RECT 49.235 96.945 50.545 97.095 ;
      RECT 49.235 97.095 50.695 97.245 ;
      RECT 49.235 97.245 50.845 97.395 ;
      RECT 49.235 97.395 50.995 97.545 ;
      RECT 49.235 97.545 51.145 97.695 ;
      RECT 49.235 97.695 51.295 97.845 ;
      RECT 49.235 97.845 51.445 97.995 ;
      RECT 49.235 97.995 51.595 98.145 ;
      RECT 49.235 98.145 51.745 98.295 ;
      RECT 49.235 98.295 51.895 98.445 ;
      RECT 49.235 98.445 52.045 98.595 ;
      RECT 49.235 98.595 52.195 98.745 ;
      RECT 49.235 98.745 52.345 98.895 ;
      RECT 49.235 98.895 52.495 99.045 ;
      RECT 49.235 99.045 52.645 99.195 ;
      RECT 49.235 99.195 52.795 99.345 ;
      RECT 49.235 99.345 52.945 99.495 ;
      RECT 49.235 99.495 53.095 99.645 ;
      RECT 49.235 99.645 53.245 99.795 ;
      RECT 49.235 99.795 53.395 99.945 ;
      RECT 49.235 99.945 53.545 100.095 ;
      RECT 49.235 100.095 53.695 100.245 ;
      RECT 49.235 100.245 53.845 100.33 ;
      RECT 49.235 164.295 53.78 164.445 ;
      RECT 49.235 164.445 53.63 164.595 ;
      RECT 49.235 164.595 53.48 164.745 ;
      RECT 49.235 164.745 53.33 164.895 ;
      RECT 49.235 164.895 53.18 165.045 ;
      RECT 49.235 165.045 53.03 165.195 ;
      RECT 49.235 165.195 52.88 165.345 ;
      RECT 49.235 165.345 52.73 165.495 ;
      RECT 49.235 165.495 52.58 165.645 ;
      RECT 49.235 165.645 52.43 165.795 ;
      RECT 49.235 165.795 52.28 165.945 ;
      RECT 49.235 165.945 52.13 166.095 ;
      RECT 49.235 166.095 51.98 166.245 ;
      RECT 49.235 166.245 51.83 166.395 ;
      RECT 49.235 166.395 51.68 166.545 ;
      RECT 49.235 166.545 51.53 166.695 ;
      RECT 49.235 166.695 51.38 166.845 ;
      RECT 49.235 166.845 51.23 166.995 ;
      RECT 49.235 166.995 51.08 167.145 ;
      RECT 49.235 167.145 50.93 167.295 ;
      RECT 49.235 167.295 50.78 167.445 ;
      RECT 49.235 167.445 50.63 167.595 ;
      RECT 49.235 167.595 50.48 167.745 ;
      RECT 49.235 167.745 50.33 167.895 ;
      RECT 49.235 167.895 50.18 168.045 ;
      RECT 49.235 168.045 50.03 168.195 ;
      RECT 49.235 168.195 49.88 168.345 ;
      RECT 49.235 168.345 49.73 168.495 ;
      RECT 49.235 168.495 49.58 168.645 ;
      RECT 49.235 168.645 49.43 168.795 ;
      RECT 49.235 168.795 49.28 168.945 ;
      RECT 49.42 84.645 75 84.795 ;
      RECT 49.57 84.795 75 84.945 ;
      RECT 49.72 84.945 75 85.095 ;
      RECT 49.87 85.095 75 85.245 ;
      RECT 50.02 85.245 75 85.395 ;
      RECT 50.17 85.395 75 85.545 ;
      RECT 50.32 85.545 75 85.695 ;
      RECT 50.47 85.695 75 85.845 ;
      RECT 50.62 85.845 75 85.995 ;
      RECT 50.77 85.995 75 86.145 ;
      RECT 50.92 86.145 75 86.295 ;
      RECT 51.07 86.295 75 86.445 ;
      RECT 51.22 86.445 75 86.595 ;
      RECT 51.37 86.595 75 86.745 ;
      RECT 51.42 86.745 75 86.795 ;
      RECT 51.57 88.21 75 88.36 ;
      RECT 51.72 88.36 75 88.51 ;
      RECT 51.87 88.51 75 88.66 ;
      RECT 52.02 88.66 75 88.81 ;
      RECT 52.17 88.81 75 88.96 ;
      RECT 52.32 88.96 75 89.11 ;
      RECT 52.47 89.11 75 89.26 ;
      RECT 52.62 89.26 75 89.41 ;
      RECT 52.77 89.41 75 89.56 ;
      RECT 52.92 89.56 75 89.71 ;
      RECT 53.07 89.71 75 89.86 ;
      RECT 53.22 89.86 75 90.01 ;
      RECT 53.37 90.01 75 90.16 ;
      RECT 53.52 90.16 75 90.31 ;
      RECT 53.67 90.31 75 90.46 ;
      RECT 53.82 90.46 75 90.61 ;
      RECT 53.97 90.61 75 90.76 ;
      RECT 54.12 90.76 75 90.91 ;
      RECT 54.27 90.91 75 91.06 ;
      RECT 54.42 91.06 75 91.21 ;
      RECT 54.57 91.21 75 91.36 ;
      RECT 54.72 91.36 75 91.51 ;
      RECT 54.87 91.51 75 91.66 ;
      RECT 55.02 91.66 75 91.81 ;
      RECT 55.17 91.81 75 91.96 ;
      RECT 55.32 91.96 75 92.11 ;
      RECT 55.47 92.11 75 92.26 ;
      RECT 55.62 92.26 75 92.41 ;
      RECT 55.77 92.41 75 92.56 ;
      RECT 55.92 92.56 75 92.71 ;
      RECT 56.07 92.71 75 92.86 ;
      RECT 32.545 86.165 33.655 86.315 ;
      RECT 32.545 86.315 33.555 86.415 ;
      RECT 33.02 84.38 33.63 84.53 ;
      RECT 32.87 84.53 33.78 84.68 ;
      RECT 32.72 84.68 33.93 84.83 ;
      RECT 32.57 84.83 34.08 84.855 ;
      RECT 34.15 163.97 42.285 164.12 ;
      RECT 34.3 164.12 42.135 164.27 ;
      RECT 34.45 164.27 41.985 164.42 ;
      RECT 34.6 164.42 41.835 164.57 ;
      RECT 34.75 164.57 41.685 164.72 ;
      RECT 34.9 164.72 41.535 164.87 ;
      RECT 35.05 164.87 41.385 165.02 ;
      RECT 35.2 165.02 41.235 165.17 ;
      RECT 35.35 165.17 41.085 165.32 ;
      RECT 35.5 165.32 40.935 165.47 ;
      RECT 35.65 165.47 40.785 165.62 ;
      RECT 35.8 165.62 40.635 165.77 ;
      RECT 35.95 165.77 40.485 165.92 ;
      RECT 36.1 165.92 40.335 166.07 ;
      RECT 36.25 166.07 40.185 166.22 ;
      RECT 36.4 166.22 40.035 166.37 ;
      RECT 36.55 166.37 39.885 166.52 ;
      RECT 36.7 166.52 39.735 166.67 ;
      RECT 36.85 166.67 39.585 166.82 ;
      RECT 37.0 166.82 39.435 166.97 ;
      RECT 37.15 166.97 39.285 167.12 ;
      RECT 37.3 167.12 39.135 167.27 ;
      RECT 37.325 167.27 39.11 167.295 ;
      RECT 37.43 70.94 75 71.09 ;
      RECT 37.58 71.09 75 71.24 ;
      RECT 37.73 71.24 75 71.39 ;
      RECT 37.88 71.39 75 71.54 ;
      RECT 38.03 71.54 75 71.69 ;
      RECT 38.18 71.69 75 71.84 ;
      RECT 38.33 71.84 75 71.99 ;
      RECT 38.48 71.99 75 72.14 ;
      RECT 38.63 72.14 75 72.29 ;
      RECT 38.78 72.29 75 72.44 ;
      RECT 38.93 72.44 75 72.59 ;
      RECT 39.08 72.59 75 72.74 ;
      RECT 39.23 72.74 75 72.89 ;
      RECT 39.38 72.89 75 73.04 ;
      RECT 39.53 73.04 75 73.19 ;
      RECT 39.68 73.19 75 73.34 ;
      RECT 39.83 73.34 75 73.49 ;
      RECT 39.98 73.49 75 73.64 ;
      RECT 40.13 73.64 75 73.79 ;
      RECT 40.28 73.79 75 73.94 ;
      RECT 40.43 73.94 75 74.09 ;
      RECT 40.58 74.09 75 74.24 ;
      RECT 40.68 74.24 75 74.34 ;
      RECT 37.325 167.295 38.96 167.445 ;
      RECT 37.325 167.445 38.81 167.595 ;
      RECT 37.325 167.595 38.66 167.745 ;
      RECT 37.325 167.745 38.51 167.895 ;
      RECT 37.325 167.895 38.36 168.045 ;
      RECT 37.325 168.045 38.21 168.195 ;
      RECT 37.325 168.195 38.06 168.345 ;
      RECT 37.325 168.345 37.91 168.495 ;
      RECT 37.325 168.495 37.76 168.645 ;
      RECT 37.325 168.645 37.61 168.795 ;
      RECT 37.325 168.795 37.46 168.945 ;
      RECT 39.935 87.195 41.21 87.345 ;
      RECT 40.085 87.345 41.21 87.495 ;
      RECT 40.2 87.495 41.21 87.61 ;
      RECT 40.26 84.38 40.735 84.53 ;
      RECT 40.11 84.53 40.885 84.68 ;
      RECT 39.96 84.68 41.035 84.83 ;
      RECT 39.81 84.83 41.185 84.855 ;
      RECT 40.35 87.61 41.21 87.76 ;
      RECT 40.5 87.76 41.36 87.91 ;
      RECT 40.65 87.91 41.51 88.06 ;
      RECT 40.8 88.06 41.66 88.21 ;
      RECT 40.95 88.21 41.81 88.36 ;
      RECT 41.1 88.36 41.96 88.51 ;
      RECT 41.25 88.51 42.11 88.66 ;
      RECT 41.4 88.66 42.26 88.81 ;
      RECT 41.55 88.81 42.41 88.96 ;
      RECT 41.7 88.96 42.56 89.11 ;
      RECT 41.85 89.11 42.71 89.26 ;
      RECT 42.0 89.26 42.86 89.41 ;
      RECT 42.15 89.41 43.01 89.56 ;
      RECT 42.3 89.56 43.16 89.71 ;
      RECT 42.45 89.71 43.31 89.86 ;
      RECT 42.6 89.86 43.46 90.01 ;
      RECT 42.75 90.01 43.61 90.16 ;
      RECT 42.9 90.16 43.76 90.31 ;
      RECT 43.05 90.31 43.91 90.46 ;
      RECT 43.2 90.46 44.06 90.61 ;
      RECT 43.35 90.61 44.21 90.76 ;
      RECT 43.5 90.76 44.36 90.91 ;
      RECT 43.65 90.91 44.51 91.06 ;
      RECT 43.8 91.06 44.66 91.21 ;
      RECT 43.95 91.21 44.81 91.36 ;
      RECT 44.1 91.36 44.96 91.51 ;
      RECT 44.25 91.51 45.11 91.66 ;
      RECT 44.4 91.66 45.26 91.81 ;
      RECT 44.55 91.81 45.41 91.96 ;
      RECT 44.7 91.96 45.56 92.11 ;
      RECT 44.85 92.11 45.71 92.26 ;
      RECT 45.0 92.26 45.86 92.41 ;
      RECT 45.15 92.41 46.01 92.56 ;
      RECT 45.3 92.56 46.16 92.71 ;
      RECT 45.45 92.71 46.31 92.86 ;
      RECT 45.6 92.86 46.46 93.01 ;
      RECT 45.75 93.01 46.61 93.16 ;
      RECT 45.9 93.16 46.76 93.31 ;
      RECT 46.05 93.31 46.91 93.46 ;
      RECT 46.2 93.46 47.06 93.61 ;
      RECT 46.35 93.61 47.21 93.76 ;
      RECT 46.5 93.76 47.36 93.91 ;
      RECT 46.65 93.91 47.51 94.06 ;
      RECT 46.8 94.06 47.66 94.21 ;
      RECT 46.95 94.21 47.81 94.36 ;
      RECT 47.1 94.36 47.96 94.51 ;
      RECT 47.25 94.51 48.11 94.66 ;
      RECT 47.4 94.66 48.26 94.81 ;
      RECT 47.55 94.81 48.41 94.96 ;
      RECT 47.7 94.96 48.56 95.11 ;
      RECT 47.85 95.11 48.71 95.26 ;
      RECT 48.0 95.26 48.86 95.41 ;
      RECT 48.15 95.41 49.01 95.56 ;
      RECT 48.3 95.56 49.16 95.71 ;
      RECT 24.855 169.635 25.635 169.785 ;
      RECT 25.005 169.785 25.635 169.935 ;
      RECT 25.155 169.935 25.635 170.085 ;
      RECT 25.305 170.085 25.635 170.235 ;
      RECT 25.455 170.235 25.635 170.385 ;
      RECT 25.605 170.385 25.635 170.535 ;
      RECT 24.625 94.335 25.635 94.485 ;
      RECT 24.475 94.485 25.635 94.635 ;
      RECT 24.325 94.635 25.635 94.785 ;
      RECT 24.175 94.785 25.635 94.935 ;
      RECT 24.025 94.935 25.635 95.085 ;
      RECT 23.875 95.085 25.635 95.235 ;
      RECT 23.725 95.235 25.635 95.385 ;
      RECT 23.575 95.385 25.635 95.535 ;
      RECT 23.425 95.535 25.635 95.685 ;
      RECT 23.275 95.685 25.635 95.835 ;
      RECT 23.125 95.835 25.635 95.985 ;
      RECT 22.975 95.985 25.635 96.135 ;
      RECT 22.825 96.135 25.635 96.285 ;
      RECT 22.675 96.285 25.635 96.435 ;
      RECT 22.525 96.435 25.635 96.585 ;
      RECT 22.375 96.585 25.635 96.735 ;
      RECT 22.225 96.735 25.635 96.885 ;
      RECT 22.075 96.885 25.635 96.955 ;
      RECT 32.545 86.415 33.405 86.565 ;
      RECT 32.395 86.565 33.255 86.715 ;
      RECT 32.245 86.715 33.105 86.865 ;
      RECT 32.095 86.865 32.955 87.015 ;
      RECT 31.945 87.015 32.805 87.165 ;
      RECT 31.795 87.165 32.655 87.315 ;
      RECT 31.645 87.315 32.505 87.465 ;
      RECT 31.495 87.465 32.355 87.615 ;
      RECT 31.345 87.615 32.205 87.765 ;
      RECT 31.195 87.765 32.055 87.915 ;
      RECT 31.045 87.915 31.905 88.065 ;
      RECT 30.895 88.065 31.755 88.215 ;
      RECT 30.745 88.215 31.605 88.365 ;
      RECT 30.595 88.365 31.455 88.515 ;
      RECT 30.445 88.515 31.305 88.665 ;
      RECT 30.295 88.665 31.155 88.815 ;
      RECT 30.145 88.815 31.005 88.965 ;
      RECT 29.995 88.965 30.855 89.115 ;
      RECT 29.845 89.115 30.705 89.265 ;
      RECT 29.695 89.265 30.555 89.415 ;
      RECT 29.545 89.415 30.405 89.565 ;
      RECT 29.395 89.565 30.255 89.715 ;
      RECT 29.245 89.715 30.105 89.865 ;
      RECT 29.095 89.865 29.955 90.015 ;
      RECT 28.945 90.015 29.805 90.165 ;
      RECT 28.795 90.165 29.655 90.315 ;
      RECT 28.645 90.315 29.505 90.465 ;
      RECT 28.495 90.465 29.355 90.615 ;
      RECT 28.345 90.615 29.205 90.765 ;
      RECT 28.195 90.765 29.055 90.915 ;
      RECT 28.045 90.915 28.905 91.065 ;
      RECT 27.895 91.065 28.755 91.215 ;
      RECT 27.745 91.215 28.605 91.365 ;
      RECT 27.595 91.365 28.455 91.515 ;
      RECT 27.445 91.515 28.305 91.665 ;
      RECT 27.295 91.665 28.155 91.815 ;
      RECT 27.145 91.815 28.005 91.965 ;
      RECT 26.995 91.965 27.855 92.115 ;
      RECT 26.845 92.115 27.705 92.265 ;
      RECT 26.695 92.265 27.555 92.415 ;
      RECT 26.545 92.415 27.405 92.565 ;
      RECT 26.395 92.565 27.255 92.715 ;
      RECT 26.245 92.715 27.105 92.865 ;
      RECT 26.095 92.865 26.955 93.015 ;
      RECT 25.945 93.015 26.805 93.165 ;
      RECT 25.795 93.165 26.655 93.315 ;
      RECT 25.645 93.315 26.505 93.465 ;
      RECT 25.495 93.465 26.355 93.615 ;
      RECT 25.345 93.615 26.205 93.765 ;
      RECT 25.195 93.765 26.055 93.915 ;
      RECT 25.045 93.915 25.905 94.065 ;
      RECT 24.895 94.065 25.755 94.215 ;
      RECT 24.745 94.215 25.635 94.335 ;
      RECT 35.215 90.775 37.63 90.925 ;
      RECT 35.065 90.925 37.78 91.075 ;
      RECT 34.915 91.075 37.93 91.225 ;
      RECT 34.765 91.225 38.08 91.375 ;
      RECT 34.615 91.375 38.23 91.525 ;
      RECT 34.465 91.525 38.38 91.675 ;
      RECT 34.315 91.675 38.53 91.825 ;
      RECT 34.165 91.825 38.68 91.975 ;
      RECT 34.015 91.975 38.83 92.125 ;
      RECT 33.865 92.125 38.98 92.275 ;
      RECT 33.715 92.275 39.13 92.425 ;
      RECT 33.565 92.425 39.28 92.575 ;
      RECT 33.415 92.575 39.43 92.725 ;
      RECT 33.265 92.725 39.58 92.875 ;
      RECT 33.115 92.875 39.73 93.025 ;
      RECT 32.965 93.025 39.88 93.175 ;
      RECT 32.815 93.175 40.03 93.325 ;
      RECT 32.665 93.325 40.18 93.475 ;
      RECT 32.515 93.475 40.33 93.555 ;
      RECT 32.435 93.555 40.41 93.705 ;
      RECT 32.435 93.705 40.56 93.855 ;
      RECT 32.435 93.855 40.71 94.005 ;
      RECT 32.435 94.005 40.86 94.155 ;
      RECT 32.435 94.155 41.01 94.305 ;
      RECT 32.435 94.305 41.16 94.455 ;
      RECT 32.435 94.455 41.31 94.605 ;
      RECT 32.435 94.605 41.46 94.755 ;
      RECT 32.435 94.755 41.61 94.905 ;
      RECT 32.435 94.905 41.76 95.055 ;
      RECT 32.435 95.055 41.91 95.205 ;
      RECT 32.435 95.205 42.06 95.355 ;
      RECT 32.435 95.355 42.21 95.505 ;
      RECT 32.435 95.505 42.36 95.58 ;
      RECT 32.585 162.405 42.435 162.555 ;
      RECT 32.735 162.555 42.435 162.705 ;
      RECT 32.885 162.705 42.435 162.855 ;
      RECT 33.035 162.855 42.435 163.005 ;
      RECT 33.185 163.005 42.435 163.155 ;
      RECT 33.335 163.155 42.435 163.305 ;
      RECT 33.485 163.305 42.435 163.455 ;
      RECT 33.635 163.455 42.435 163.605 ;
      RECT 33.785 163.605 42.435 163.755 ;
      RECT 33.935 163.755 42.435 163.905 ;
      RECT 34.0 163.905 42.435 163.97 ;
      RECT 32.545 85.865 33.955 86.015 ;
      RECT 32.545 86.015 33.805 86.165 ;
      RECT 32.545 84.855 34.105 85.865 ;
      RECT 39.785 84.855 41.21 87.195 ;
      RECT 0 0 24.64 3.005 ;
      RECT 0 3.005 3.005 82.335 ;
      RECT 0 84.485 3.0 85.9 ;
      RECT 15.205 194.995 60.73 198 ;
      RECT 15.205 189.915 60.73 192.92 ;
      RECT 20.45 84.485 23.45 84.655 ;
      RECT 21.355 79.33 25.6 82.335 ;
      RECT 21.635 3.005 24.64 24.785 ;
      RECT 21.64 24.785 25.6 27.79 ;
      RECT 22.005 96.955 25.635 166.935 ;
      RECT 22.595 27.79 25.6 79.33 ;
      RECT 32.435 95.58 42.435 162.405 ;
      RECT 37.28 0 37.98 69.89 ;
      RECT 37.28 69.89 52.66 70.94 ;
      RECT 49.235 100.33 53.93 164.295 ;
      RECT 49.27 81.64 53.515 84.645 ;
      RECT 49.27 76.65 52.275 81.64 ;
      RECT 49.655 3.005 52.66 69.89 ;
      RECT 49.655 70.94 52.66 74.34 ;
      RECT 49.655 0 75 3.005 ;
      RECT 51.42 86.795 54.42 86.965 ;
      RECT 71.995 76.65 75 84.645 ;
      RECT 71.995 3.005 75 74.34 ;
      RECT 72.0 86.795 75 88.21 ;
      RECT 3.0 83.24 20.45 84.655 ;
      RECT 3.0 27.785 22.595 81.09 ;
      RECT 3.0 3.002 21.64 27.785 ;
      RECT 0 94.145 15.205 198 ;
      RECT 3.0 92.9 12.205 192.915 ;
      RECT 52.27 75.405 72.0 83.4 ;
      RECT 54.42 85.55 72.0 86.965 ;
      RECT 3.0 192.915 72.0 195.0 ;
      RECT 60.73 97.52 75 198 ;
      RECT 63.73 96.275 72.0 192.915 ;
      RECT 52.655 3.0 72.0 72.89 ;
      RECT 0 85.9 23.3 86.05 ;
      RECT 0 86.05 23.15 86.2 ;
      RECT 0 86.2 23.0 86.35 ;
      RECT 0 86.35 22.85 86.5 ;
      RECT 0 86.5 22.7 86.65 ;
      RECT 0 86.65 22.55 86.8 ;
      RECT 0 86.8 22.4 86.95 ;
      RECT 0 86.95 22.25 87.1 ;
      RECT 0 87.1 22.1 87.25 ;
      RECT 0 87.25 21.95 87.4 ;
      RECT 0 87.4 21.8 87.55 ;
      RECT 0 87.55 21.65 87.7 ;
      RECT 0 87.7 21.5 87.85 ;
      RECT 0 87.85 21.35 88 ;
      RECT 0 88 21.2 88.15 ;
      RECT 0 88.15 21.05 88.3 ;
      RECT 0 88.3 20.9 88.45 ;
      RECT 0 88.45 20.75 88.6 ;
      RECT 0 88.6 20.6 88.75 ;
      RECT 0 88.75 20.45 88.9 ;
      RECT 0 88.9 20.3 89.05 ;
      RECT 0 89.05 20.15 89.2 ;
      RECT 0 89.2 20.0 89.35 ;
      RECT 0 89.35 19.85 89.5 ;
      RECT 0 89.5 19.7 89.65 ;
      RECT 0 89.65 19.55 89.8 ;
      RECT 0 89.8 19.4 89.95 ;
      RECT 0 89.95 19.25 90.1 ;
      RECT 0 90.1 19.1 90.25 ;
      RECT 0 90.25 18.95 90.4 ;
      RECT 0 90.4 18.8 90.55 ;
      RECT 0 90.55 18.65 90.7 ;
      RECT 0 90.7 18.5 90.85 ;
      RECT 0 90.85 18.35 91 ;
      RECT 0 91 18.2 91.15 ;
      RECT 0 91.15 18.05 91.3 ;
      RECT 0 91.3 17.9 91.45 ;
      RECT 0 91.45 17.75 91.6 ;
      RECT 0 91.6 17.6 91.75 ;
      RECT 0 91.75 17.45 91.9 ;
      RECT 0 91.9 17.3 92.05 ;
      RECT 0 92.05 17.15 92.2 ;
      RECT 0 92.2 17.0 92.35 ;
      RECT 0 92.35 16.85 92.5 ;
      RECT 0 92.5 16.7 92.65 ;
      RECT 0 92.65 16.55 92.8 ;
      RECT 0 92.8 16.4 92.95 ;
      RECT 0 92.95 16.25 93.1 ;
      RECT 0 93.1 16.1 93.25 ;
      RECT 0 93.25 15.95 93.4 ;
      RECT 0 93.4 15.8 93.55 ;
      RECT 0 93.55 15.65 93.7 ;
      RECT 0 93.7 15.5 93.85 ;
      RECT 0 93.85 15.35 94 ;
      RECT 0 94 15.205 94.145 ;
      RECT 0 82.335 25.45 82.485 ;
      RECT 0 82.485 25.3 82.635 ;
      RECT 0 82.635 25.15 82.785 ;
      RECT 0 82.785 25.0 82.935 ;
      RECT 0 82.935 24.85 83.085 ;
      RECT 0 83.085 24.7 83.235 ;
      RECT 0 83.235 24.55 83.385 ;
      RECT 0 83.385 24.4 83.535 ;
      RECT 0 83.535 24.25 83.685 ;
      RECT 0 83.685 24.1 83.835 ;
      RECT 0 83.835 23.95 83.985 ;
      RECT 0 83.985 23.8 84.135 ;
      RECT 0 84.135 23.65 84.285 ;
      RECT 0 84.285 23.5 84.435 ;
      RECT 0 84.435 23.45 84.485 ;
      RECT 22.155 166.935 25.635 167.085 ;
      RECT 22.305 167.085 25.635 167.235 ;
      RECT 22.455 167.235 25.635 167.385 ;
      RECT 22.605 167.385 25.635 167.535 ;
      RECT 22.755 167.535 25.635 167.685 ;
      RECT 22.905 167.685 25.635 167.835 ;
      RECT 23.055 167.835 25.635 167.985 ;
      RECT 23.205 167.985 25.635 168.135 ;
      RECT 23.355 168.135 25.635 168.285 ;
      RECT 23.505 168.285 25.635 168.435 ;
      RECT 23.655 168.435 25.635 168.585 ;
      RECT 23.805 168.585 25.635 168.735 ;
      RECT 23.955 168.735 25.635 168.885 ;
      RECT 24.105 168.885 25.635 169.035 ;
      RECT 24.255 169.035 25.635 169.185 ;
      RECT 24.405 169.185 25.635 169.335 ;
      RECT 24.555 169.335 25.635 169.485 ;
      RECT 24.705 169.485 25.635 169.635 ;
    LAYER met5 ;
      RECT 0 0 75 198 ;
    LAYER met4 ;
      RECT 0 0 75 198 ;
  END
END sky130_fd_io__top_lvc_b2b
  
END LIBRARY
