# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_gpiov2
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_gpiov2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  80.00000 BY  200.0000 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.760000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.465000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430000 0.000000 62.690000 1.305000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865000 0.000000 46.195000 36.805000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.750000 0.000000 31.010000 2.265000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.855000 0.000000 50.115000 0.545000 ;
    END
  END DM[0]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.835000 0.000000 67.095000 1.195000 ;
    END
  END DM[1]
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490000 0.000000 28.750000 4.070000 ;
    END
  END DM[2]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.460000 0.000000 35.720000 1.550000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390000 0.000000 38.650000 3.090000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.755000 0.000000 13.015000 5.350000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580000 0.000000 78.910000 184.775000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.310000 0.000000 16.570000 2.320000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815000 0.000000 32.075000 3.340000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600000 0.000000 26.860000 2.705000 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420000 0.000000 5.650000 4.475000 ;
    END
  END IB_MODE_SEL
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240000 0.000000 79.570000 189.560000 ;
    END
  END IN
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245000 0.000000 45.505000 5.090000 ;
    END
  END INP_DIS
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400000 0.000000 1.020000 178.485000 ;
    END
  END IN_H
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375000 0.000000 3.605000 4.475000 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355000 0.000000 22.615000 6.425000 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.100000 104.395000 73.800000 167.010000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280000 0.000000 76.920000 2.055000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275000 0.000000 68.925000 2.270000 ;
    END
    PORT
      LAYER met2 ;
        RECT 68.405000 0.105000 68.415000 0.115000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000000 106.585000 12.500000 118.955000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.515000 118.955000 8.570000 120.010000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.665000 118.955000 12.500000 119.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.815000 119.105000 12.500000 119.255000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.830000 106.210000 8.205000 106.585000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.850000 106.565000 12.500000 106.585000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.965000 119.255000 12.500000 119.405000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.000000 106.415000 12.500000 106.565000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.115000 119.405000 12.500000 119.555000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.205000 105.030000 9.385000 106.210000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.265000 119.555000 12.500000 119.705000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.300000 106.115000 12.500000 106.265000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.415000 119.705000 12.500000 119.855000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.450000 105.965000 12.500000 106.115000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.570000 120.010000 9.800000 121.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.600000 105.815000 12.500000 105.965000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.715000 120.005000 12.500000 120.155000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.750000 105.665000 12.500000 105.815000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.865000 120.155000 12.500000 120.305000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.900000 105.515000 12.500000 105.665000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.015000 120.305000 12.500000 120.455000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.050000 105.365000 12.500000 105.515000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.165000 120.455000 12.500000 120.605000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.200000 105.215000 12.500000 105.365000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.315000 120.605000 12.500000 120.755000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.385000 104.395000 10.020000 105.030000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.465000 120.755000 12.500000 120.905000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.500000 104.915000 12.500000 105.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.615000 120.905000 12.500000 121.055000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.650000 104.765000 12.500000 104.915000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.810000 121.205000 12.500000 121.250000 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.610000 0.000000 77.870000 1.185000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.705000 0.000000 78.905000 1.215000 ;
    END
    PORT
      LAYER met2 ;
        RECT 78.800000 0.105000 78.810000 0.115000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715000 0.000000 79.915000 177.870000 ;
    END
  END TIE_LO_ESD
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130000 0.000000 6.390000 1.550000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 70.265000 8.885000 80.000000 13.535000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 76.810000 2.035000 80.000000 7.485000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 51.570000 14.935000 80.000000 18.385000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 68.030000 70.035000 80.000000 95.000000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 60.945000 64.085000 80.000000 68.535000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 47.090000 56.405000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 55.705000 41.585000 80.000000 46.235000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.530000 25.835000 80.000000 30.485000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 71.575000 58.235000 80.000000 62.685000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.850000 31.885000 80.000000 35.335000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT 0.000000 0.230000 80.000000 199.705000 ;
    LAYER met1 ;
      RECT  0.000000 0.260000 62.150000   1.585000 ;
      RECT  0.000000 1.585000 80.000000 200.000000 ;
      RECT 62.970000 0.260000 80.000000   1.585000 ;
    LAYER met2 ;
      RECT  0.210000   0.250000  3.095000   4.755000 ;
      RECT  0.210000   4.755000 12.475000   5.630000 ;
      RECT  0.210000   5.630000 22.075000   6.705000 ;
      RECT  0.210000   6.705000 79.435000 178.150000 ;
      RECT  0.210000 178.150000 79.915000 200.000000 ;
      RECT  3.885000   0.250000  5.140000   4.755000 ;
      RECT  5.930000   1.830000 12.475000   4.755000 ;
      RECT  6.670000   0.250000 12.475000   1.830000 ;
      RECT 13.295000   0.250000 16.030000   2.600000 ;
      RECT 13.295000   2.600000 22.075000   5.630000 ;
      RECT 16.850000   0.250000 22.075000   2.600000 ;
      RECT 22.895000   0.250000 26.320000   2.985000 ;
      RECT 22.895000   2.985000 28.210000   4.350000 ;
      RECT 22.895000   4.350000 44.965000   5.370000 ;
      RECT 22.895000   5.370000 79.435000   6.705000 ;
      RECT 27.140000   0.250000 28.210000   2.985000 ;
      RECT 29.030000   0.250000 30.470000   2.545000 ;
      RECT 29.030000   2.545000 31.535000   3.620000 ;
      RECT 29.030000   3.620000 44.965000   4.350000 ;
      RECT 31.290000   0.250000 31.535000   2.545000 ;
      RECT 32.355000   0.250000 35.180000   1.830000 ;
      RECT 32.355000   1.830000 38.110000   3.370000 ;
      RECT 32.355000   3.370000 44.965000   3.620000 ;
      RECT 36.000000   0.250000 38.110000   1.830000 ;
      RECT 38.930000   0.250000 44.965000   3.370000 ;
      RECT 45.785000   0.250000 49.575000   0.825000 ;
      RECT 45.785000   0.825000 66.555000   1.475000 ;
      RECT 45.785000   1.475000 67.995000   2.550000 ;
      RECT 45.785000   2.550000 79.435000   5.370000 ;
      RECT 50.395000   0.250000 66.555000   0.825000 ;
      RECT 67.375000   0.250000 67.995000   1.475000 ;
      RECT 69.205000   0.250000 76.000000   2.335000 ;
      RECT 69.205000   2.335000 79.435000   2.550000 ;
      RECT 77.200000   0.250000 77.330000   1.465000 ;
      RECT 77.200000   1.465000 78.425000   1.495000 ;
      RECT 77.200000   1.495000 79.435000   2.335000 ;
      RECT 78.150000   0.250000 78.425000   1.465000 ;
      RECT 79.185000   0.250000 79.435000   1.495000 ;
    LAYER met3 ;
      RECT  0.400000 178.885000 78.180000 185.175000 ;
      RECT  0.400000 185.175000 78.840000 189.960000 ;
      RECT  0.400000 189.960000 79.570000 200.000000 ;
      RECT  1.420000   0.000000 45.465000  37.205000 ;
      RECT  1.420000  37.205000 78.180000 178.885000 ;
      RECT 46.595000   0.000000 78.180000  37.205000 ;
    LAYER met4 ;
      RECT  0.000000   0.535000 80.000000   1.635000 ;
      RECT  0.000000   1.635000 76.410000   7.885000 ;
      RECT  0.000000   7.885000 80.000000   8.485000 ;
      RECT  0.000000   8.485000 69.865000  13.935000 ;
      RECT  0.000000  13.935000 80.000000  14.535000 ;
      RECT  0.000000  14.535000 51.170000  18.785000 ;
      RECT  0.000000  18.785000 80.000000  25.435000 ;
      RECT  0.000000  25.435000 21.130000  30.885000 ;
      RECT  0.000000  30.885000 80.000000  31.485000 ;
      RECT  0.000000  31.485000 23.450000  35.735000 ;
      RECT  0.000000  35.735000 80.000000  41.185000 ;
      RECT  0.000000  41.185000 55.305000  46.635000 ;
      RECT  0.000000  46.635000 80.000000  47.965000 ;
      RECT  0.000000  47.965000 54.065000  51.745000 ;
      RECT  0.000000  51.745000 80.000000  52.725000 ;
      RECT  0.000000  52.725000 38.360000  56.505000 ;
      RECT  0.000000  56.505000 46.690000  57.135000 ;
      RECT  0.000000  57.135000 80.000000  57.835000 ;
      RECT  0.000000  57.835000 71.175000  63.085000 ;
      RECT  0.000000  63.085000 80.000000  63.685000 ;
      RECT  0.000000  63.685000 60.545000  68.935000 ;
      RECT  0.000000  68.935000 80.000000  69.635000 ;
      RECT  0.000000  69.635000 67.630000  95.400000 ;
      RECT  0.000000  95.400000 80.000000 103.995000 ;
      RECT  0.000000 103.995000  8.985000 104.630000 ;
      RECT  0.000000 104.630000  7.805000 105.810000 ;
      RECT  0.000000 105.810000  7.430000 106.185000 ;
      RECT  0.000000 106.185000  1.600000 119.355000 ;
      RECT  0.000000 119.355000  7.115000 120.410000 ;
      RECT  0.000000 120.410000  8.170000 121.640000 ;
      RECT  0.000000 121.640000  9.410000 121.650000 ;
      RECT  0.000000 121.650000 80.000000 200.000000 ;
      RECT 10.420000 103.995000 80.000000 104.365000 ;
      RECT 12.900000 104.365000 80.000000 121.650000 ;
    LAYER met5 ;
      RECT 9.800000  98.085000 75.200000 102.795000 ;
      RECT 9.800000 168.610000 75.200000 173.485000 ;
  END
END sky130_fd_io__top_gpiov2
END LIBRARY
